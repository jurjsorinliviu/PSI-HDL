* ngspice behavioral subcircuit (B-sources)
* Generated from model: PsiNN_burgers
.subckt psi_nn_psinn_burgers in0 in1 out0 vdd vss

* Activation (fallback-friendly): use tanh() if supported by ngspice, else replace with rational approx
.func tanh_psi(x) { tanh(x) }

B_u1p_0 u1p_0 0 V = tanh_psi(8.668856620789e-01 + -3.981690406799e-01*V(in0) + -1.969884634018e-01*V(in1))
B_u1m_0 u1m_0 0 V = tanh_psi(8.668856620789e-01 + -3.981690406799e-01*V(in0) + (-1)*(-1.969884634018e-01*V(in1)))
B_u1p_1 u1p_1 0 V = tanh_psi(6.342871189117e-01 + -8.205217123032e-01*V(in0) + 7.848736047745e-01*V(in1))
B_u1m_1 u1m_1 0 V = tanh_psi(6.342871189117e-01 + -8.205217123032e-01*V(in0) + (-1)*(7.848736047745e-01*V(in1)))
B_u1p_2 u1p_2 0 V = tanh_psi(9.264670610428e-01 + -3.798186779022e-02*V(in0) + -8.483624458313e-02*V(in1))
B_u1m_2 u1m_2 0 V = tanh_psi(9.264670610428e-01 + -3.798186779022e-02*V(in0) + (-1)*(-8.483624458313e-02*V(in1)))
B_u1p_3 u1p_3 0 V = tanh_psi(3.785117864609e-01 + -8.562246561050e-01*V(in0) + 7.593704462051e-01*V(in1))
B_u1m_3 u1m_3 0 V = tanh_psi(3.785117864609e-01 + -8.562246561050e-01*V(in0) + (-1)*(7.593704462051e-01*V(in1)))
B_u1p_4 u1p_4 0 V = tanh_psi(-6.512863636017e-01 + 9.649646282196e-02*V(in0) + -4.379376173019e-01*V(in1))
B_u1m_4 u1m_4 0 V = tanh_psi(-6.512863636017e-01 + 9.649646282196e-02*V(in0) + (-1)*(-4.379376173019e-01*V(in1)))
B_u1p_5 u1p_5 0 V = tanh_psi(1.098680496216e-02 + -2.397497892380e-01*V(in0) + 4.065411090851e-01*V(in1))
B_u1m_5 u1m_5 0 V = tanh_psi(1.098680496216e-02 + -2.397497892380e-01*V(in0) + (-1)*(4.065411090851e-01*V(in1)))
B_u1p_6 u1p_6 0 V = tanh_psi(5.707535743713e-01 + -6.759240627289e-01*V(in0) + -8.787122964859e-01*V(in1))
B_u1m_6 u1m_6 0 V = tanh_psi(5.707535743713e-01 + -6.759240627289e-01*V(in0) + (-1)*(-8.787122964859e-01*V(in1)))
B_u1p_7 u1p_7 0 V = tanh_psi(-9.706660509109e-01 + -9.442222118378e-02*V(in0) + -3.238424062729e-01*V(in1))
B_u1m_7 u1m_7 0 V = tanh_psi(-9.706660509109e-01 + -9.442222118378e-02*V(in0) + (-1)*(-3.238424062729e-01*V(in1)))
B_u1p_8 u1p_8 0 V = tanh_psi(-6.885164976120e-01 + 3.249348402023e-01*V(in0) + 9.765121936798e-01*V(in1))
B_u1m_8 u1m_8 0 V = tanh_psi(-6.885164976120e-01 + 3.249348402023e-01*V(in0) + (-1)*(9.765121936798e-01*V(in1)))
B_u1p_9 u1p_9 0 V = tanh_psi(-8.247464895248e-01 + -2.036794424057e-01*V(in0) + 9.787846803665e-01*V(in1))
B_u1m_9 u1m_9 0 V = tanh_psi(-8.247464895248e-01 + -2.036794424057e-01*V(in0) + (-1)*(9.787846803665e-01*V(in1)))
B_u1p_10 u1p_10 0 V = tanh_psi(2.567453384399e-01 + 4.302449226379e-01*V(in0) + -8.005249500275e-02*V(in1))
B_u1m_10 u1m_10 0 V = tanh_psi(2.567453384399e-01 + 4.302449226379e-01*V(in0) + (-1)*(-8.005249500275e-02*V(in1)))
B_u1p_11 u1p_11 0 V = tanh_psi(8.087372779846e-01 + 4.807125329971e-01*V(in0) + -1.358202695847e-01*V(in1))
B_u1m_11 u1m_11 0 V = tanh_psi(8.087372779846e-01 + 4.807125329971e-01*V(in0) + (-1)*(-1.358202695847e-01*V(in1)))
B_u1p_12 u1p_12 0 V = tanh_psi(-5.975322723389e-01 + 6.096847057343e-01*V(in0) + 5.500133037567e-01*V(in1))
B_u1m_12 u1m_12 0 V = tanh_psi(-5.975322723389e-01 + 6.096847057343e-01*V(in0) + (-1)*(5.500133037567e-01*V(in1)))
B_u1p_13 u1p_13 0 V = tanh_psi(-3.085759878159e-01 + 4.325067996979e-02*V(in0) + -4.672693014145e-01*V(in1))
B_u1m_13 u1m_13 0 V = tanh_psi(-3.085759878159e-01 + 4.325067996979e-02*V(in0) + (-1)*(-4.672693014145e-01*V(in1)))
B_u1p_14 u1p_14 0 V = tanh_psi(-9.933235645294e-01 + 6.558771133423e-01*V(in0) + 4.463710784912e-01*V(in1))
B_u1m_14 u1m_14 0 V = tanh_psi(-9.933235645294e-01 + 6.558771133423e-01*V(in0) + (-1)*(4.463710784912e-01*V(in1)))
B_u1p_15 u1p_15 0 V = tanh_psi(-3.185240030289e-01 + 6.553682088852e-01*V(in0) + -2.739950418472e-01*V(in1))
B_u1m_15 u1m_15 0 V = tanh_psi(-3.185240030289e-01 + 6.553682088852e-01*V(in0) + (-1)*(-2.739950418472e-01*V(in1)))
B_u1p_16 u1p_16 0 V = tanh_psi(-9.608575105667e-01 + -8.734289407730e-01*V(in0) + 9.083031415939e-01*V(in1))
B_u1m_16 u1m_16 0 V = tanh_psi(-9.608575105667e-01 + -8.734289407730e-01*V(in0) + (-1)*(9.083031415939e-01*V(in1)))
B_u1p_17 u1p_17 0 V = tanh_psi(4.706679582596e-01 + 2.024590969086e-02*V(in0) + -9.608633518219e-01*V(in1))
B_u1m_17 u1m_17 0 V = tanh_psi(4.706679582596e-01 + 2.024590969086e-02*V(in0) + (-1)*(-9.608633518219e-01*V(in1)))
B_u1p_18 u1p_18 0 V = tanh_psi(-6.856670379639e-01 + -1.681953668594e-01*V(in0) + 8.587348461151e-02*V(in1))
B_u1m_18 u1m_18 0 V = tanh_psi(-6.856670379639e-01 + -1.681953668594e-01*V(in0) + (-1)*(8.587348461151e-02*V(in1)))
B_u1p_19 u1p_19 0 V = tanh_psi(-6.401425600052e-01 + 1.162674427032e-01*V(in0) + -7.768144607544e-01*V(in1))
B_u1m_19 u1m_19 0 V = tanh_psi(-6.401425600052e-01 + 1.162674427032e-01*V(in0) + (-1)*(-7.768144607544e-01*V(in1)))
B_u2a_0 u2a_0 0 V = tanh_psi(5.034162104130e-02 + 2.128101587296e-01*V(u1p_0) + 1.705591678619e-01*V(u1p_1) + -1.660106480122e-01*V(u1p_2)
+ + 1.452274620533e-01*V(u1p_3) + -1.385001838207e-01*V(u1p_4) + -6.884902715683e-03*V(u1p_5) + 3.886032104492e-02*V(u1p_6)
+ + 1.961986124516e-01*V(u1p_7) + -1.448850780725e-01*V(u1p_8) + -4.922452569008e-02*V(u1p_9) + -1.904224157333e-01*V(u1p_10)
+ + -2.225336730480e-01*V(u1p_11) + -1.471883356571e-01*V(u1p_12) + -1.588267832994e-01*V(u1p_13) + 2.093329429626e-01*V(u1p_14)
+ + 1.198337674141e-01*V(u1p_15) + -1.388807594776e-02*V(u1p_16) + -2.176393568516e-02*V(u1p_17) + 1.104081571102e-01*V(u1p_18)
+ + -1.343870609999e-01*V(u1p_19) + 5.860885977745e-02*V(u1m_0) + -1.094810664654e-02*V(u1m_1) + 8.004984259605e-02*V(u1m_2)
+ + 1.569007635117e-01*V(u1m_3) + -5.736637115479e-02*V(u1m_4) + -7.305976748466e-02*V(u1m_5) + 5.592474341393e-02*V(u1m_6)
+ + 1.369167864323e-02*V(u1m_7) + 2.166581749916e-01*V(u1m_8) + 1.534524559975e-02*V(u1m_9) + 1.774801611900e-01*V(u1m_10)
+ + -2.166749536991e-01*V(u1m_11) + 2.027099132538e-01*V(u1m_12) + 1.110502779484e-01*V(u1m_13) + 4.960280656815e-02*V(u1m_14)
+ + -7.500165700912e-02*V(u1m_15) + 1.699292659760e-01*V(u1m_16) + 7.934957742691e-03*V(u1m_17) + -1.897763013840e-01*V(u1m_18)
+ + 1.165036559105e-01*V(u1m_19))
B_u2b_0 u2b_0 0 V = tanh_psi(5.034162104130e-02 + 5.860885977745e-02*V(u1p_0) + -1.094810664654e-02*V(u1p_1) + 8.004984259605e-02*V(u1p_2)
+ + 1.569007635117e-01*V(u1p_3) + -5.736637115479e-02*V(u1p_4) + -7.305976748466e-02*V(u1p_5) + 5.592474341393e-02*V(u1p_6)
+ + 1.369167864323e-02*V(u1p_7) + 2.166581749916e-01*V(u1p_8) + 1.534524559975e-02*V(u1p_9) + 1.774801611900e-01*V(u1p_10)
+ + -2.166749536991e-01*V(u1p_11) + 2.027099132538e-01*V(u1p_12) + 1.110502779484e-01*V(u1p_13) + 4.960280656815e-02*V(u1p_14)
+ + -7.500165700912e-02*V(u1p_15) + 1.699292659760e-01*V(u1p_16) + 7.934957742691e-03*V(u1p_17) + -1.897763013840e-01*V(u1p_18)
+ + 1.165036559105e-01*V(u1p_19) + 2.128101587296e-01*V(u1m_0) + 1.705591678619e-01*V(u1m_1) + -1.660106480122e-01*V(u1m_2)
+ + 1.452274620533e-01*V(u1m_3) + -1.385001838207e-01*V(u1m_4) + -6.884902715683e-03*V(u1m_5) + 3.886032104492e-02*V(u1m_6)
+ + 1.961986124516e-01*V(u1m_7) + -1.448850780725e-01*V(u1m_8) + -4.922452569008e-02*V(u1m_9) + -1.904224157333e-01*V(u1m_10)
+ + -2.225336730480e-01*V(u1m_11) + -1.471883356571e-01*V(u1m_12) + -1.588267832994e-01*V(u1m_13) + 2.093329429626e-01*V(u1m_14)
+ + 1.198337674141e-01*V(u1m_15) + -1.388807594776e-02*V(u1m_16) + -2.176393568516e-02*V(u1m_17) + 1.104081571102e-01*V(u1m_18)
+ + -1.343870609999e-01*V(u1m_19))
B_u2c_0 u2c_0 0 V = tanh_psi(0.0 + 2.067486345768e-01*(V(u1p_0) + (-1)*V(u1m_0)) + -2.261252701283e-02*(V(u1p_1) + (-1)*V(u1m_1))
+ + -1.154354140162e-01*(V(u1p_2) + (-1)*V(u1m_2)) + 1.082925498486e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.480919122696e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 2.184172868729e-01*(V(u1p_5) + (-1)*V(u1m_5)) + -1.205638125539e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + -1.390144377947e-01*(V(u1p_7) + (-1)*V(u1m_7)) + -1.186159253120e-01*(V(u1p_8) + (-1)*V(u1m_8)) + -3.173339366913e-02*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 4.454585909843e-02*(V(u1p_10) + (-1)*V(u1m_10)) + 8.521136641502e-02*(V(u1p_11) + (-1)*V(u1m_11))
+ + -2.099081724882e-01*(V(u1p_12) + (-1)*V(u1m_12)) + 6.849381327629e-02*(V(u1p_13) + (-1)*V(u1m_13)) + 1.944413781166e-01*(V(u1p_14)
+ + (-1)*V(u1m_14)) + 9.259343147278e-03*(V(u1p_15) + (-1)*V(u1m_15)) + 7.678011059761e-02*(V(u1p_16) + (-1)*V(u1m_16))
+ + -1.182915493846e-01*(V(u1p_17) + (-1)*V(u1m_17)) + 9.840413928032e-02*(V(u1p_18) + (-1)*V(u1m_18)) + 1.524708271027e-01*(V(u1p_19)
+ + (-1)*V(u1m_19)))
B_u2a_1 u2a_1 0 V = tanh_psi(1.618932932615e-01 + -2.104981243610e-01*V(u1p_0) + 1.202766895294e-01*V(u1p_1) + 1.249209046364e-02*V(u1p_2)
+ + -1.363043189049e-01*V(u1p_3) + 1.005745828152e-01*V(u1p_4) + -3.644995391369e-02*V(u1p_5) + 9.246608614922e-02*V(u1p_6)
+ + 2.189127802849e-01*V(u1p_7) + 7.821774482727e-02*V(u1p_8) + -2.894940972328e-02*V(u1p_9) + -1.611749827862e-02*V(u1p_10)
+ + -6.432281434536e-02*V(u1p_11) + 1.924041211605e-01*V(u1p_12) + -2.111572176218e-01*V(u1p_13) + 1.340722739697e-01*V(u1p_14)
+ + 8.059597015381e-02*V(u1p_15) + -1.170441284776e-01*V(u1p_16) + 2.235240340233e-01*V(u1p_17) + -4.316478967667e-02*V(u1p_18)
+ + -8.587597310543e-02*V(u1p_19) + 1.634362041950e-01*V(u1m_0) + -1.114525273442e-01*V(u1m_1) + 2.412776648998e-02*V(u1m_2)
+ + 2.319616079330e-02*V(u1m_3) + -1.975823193789e-01*V(u1m_4) + 5.406910181046e-02*V(u1m_5) + -3.069490194321e-03*V(u1m_6)
+ + 2.022019326687e-01*V(u1m_7) + -1.026756092906e-01*V(u1m_8) + -1.936025023460e-01*V(u1m_9) + -1.079176962376e-01*V(u1m_10)
+ + 8.259499073029e-02*V(u1m_11) + -1.404038071632e-01*V(u1m_12) + -1.409964263439e-01*V(u1m_13) + -7.498334348202e-02*V(u1m_14)
+ + -1.044262647629e-01*V(u1m_15) + -1.131351590157e-01*V(u1m_16) + 1.862905025482e-01*V(u1m_17) + 1.277655065060e-01*V(u1m_18)
+ + -9.052240848541e-02*V(u1m_19))
B_u2b_1 u2b_1 0 V = tanh_psi(1.618932932615e-01 + 1.634362041950e-01*V(u1p_0) + -1.114525273442e-01*V(u1p_1) + 2.412776648998e-02*V(u1p_2)
+ + 2.319616079330e-02*V(u1p_3) + -1.975823193789e-01*V(u1p_4) + 5.406910181046e-02*V(u1p_5) + -3.069490194321e-03*V(u1p_6)
+ + 2.022019326687e-01*V(u1p_7) + -1.026756092906e-01*V(u1p_8) + -1.936025023460e-01*V(u1p_9) + -1.079176962376e-01*V(u1p_10)
+ + 8.259499073029e-02*V(u1p_11) + -1.404038071632e-01*V(u1p_12) + -1.409964263439e-01*V(u1p_13) + -7.498334348202e-02*V(u1p_14)
+ + -1.044262647629e-01*V(u1p_15) + -1.131351590157e-01*V(u1p_16) + 1.862905025482e-01*V(u1p_17) + 1.277655065060e-01*V(u1p_18)
+ + -9.052240848541e-02*V(u1p_19) + -2.104981243610e-01*V(u1m_0) + 1.202766895294e-01*V(u1m_1) + 1.249209046364e-02*V(u1m_2)
+ + -1.363043189049e-01*V(u1m_3) + 1.005745828152e-01*V(u1m_4) + -3.644995391369e-02*V(u1m_5) + 9.246608614922e-02*V(u1m_6)
+ + 2.189127802849e-01*V(u1m_7) + 7.821774482727e-02*V(u1m_8) + -2.894940972328e-02*V(u1m_9) + -1.611749827862e-02*V(u1m_10)
+ + -6.432281434536e-02*V(u1m_11) + 1.924041211605e-01*V(u1m_12) + -2.111572176218e-01*V(u1m_13) + 1.340722739697e-01*V(u1m_14)
+ + 8.059597015381e-02*V(u1m_15) + -1.170441284776e-01*V(u1m_16) + 2.235240340233e-01*V(u1m_17) + -4.316478967667e-02*V(u1m_18)
+ + -8.587597310543e-02*V(u1m_19))
B_u2c_1 u2c_1 0 V = tanh_psi(0.0 + 1.322577893734e-01*(V(u1p_0) + (-1)*V(u1m_0)) + 6.117492914200e-03*(V(u1p_1) + (-1)*V(u1m_1))
+ + 5.362692475319e-02*(V(u1p_2) + (-1)*V(u1m_2)) + 3.711703419685e-02*(V(u1p_3) + (-1)*V(u1m_3)) + 2.104170322418e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + -1.129637062550e-01*(V(u1p_5) + (-1)*V(u1m_5)) + -7.027824223042e-02*(V(u1p_6) + (-1)*V(u1m_6))
+ + 2.018493413925e-02*(V(u1p_7) + (-1)*V(u1m_7)) + -1.445212364197e-01*(V(u1p_8) + (-1)*V(u1m_8)) + -1.092550158501e-02*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -1.808278262615e-01*(V(u1p_10) + (-1)*V(u1m_10)) + 1.050741672516e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + -4.420328140259e-02*(V(u1p_12) + (-1)*V(u1m_12)) + 5.615136027336e-02*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.226402893662e-01*(V(u1p_14) + (-1)*V(u1m_14)) + 1.357417702675e-01*(V(u1p_15) + (-1)*V(u1m_15))
+ + -1.005104705691e-01*(V(u1p_16) + (-1)*V(u1m_16)) + -1.534315943718e-01*(V(u1p_17) + (-1)*V(u1m_17))
+ + -1.556794941425e-01*(V(u1p_18) + (-1)*V(u1m_18)) + -1.624975800514e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_2 u2a_2 0 V = tanh_psi(-3.378880620003e-01 + 1.407382786274e-01*V(u1p_0) + 2.002112567425e-01*V(u1p_1) + 7.116436958313e-03*V(u1p_2)
+ + 2.026466131210e-01*V(u1p_3) + -8.188287913799e-02*V(u1p_4) + 3.207176923752e-03*V(u1p_5) + -3.131516277790e-02*V(u1p_6)
+ + 1.129356324673e-01*V(u1p_7) + -1.737996488810e-01*V(u1p_8) + 1.128564178944e-01*V(u1p_9) + 8.042323589325e-02*V(u1p_10)
+ + 3.867527842522e-02*V(u1p_11) + -1.359773874283e-01*V(u1p_12) + 1.179875731468e-01*V(u1p_13) + 9.016263484955e-02*V(u1p_14)
+ + -2.096267789602e-01*V(u1p_15) + -1.058997288346e-01*V(u1p_16) + -1.962925493717e-01*V(u1p_17) + -1.598631441593e-01*V(u1p_18)
+ + 7.738000154495e-02*V(u1p_19) + 1.110349297523e-01*V(u1m_0) + 3.986474871635e-02*V(u1m_1) + 2.204366326332e-01*V(u1m_2)
+ + 1.056722402573e-01*V(u1m_3) + -1.978406906128e-01*V(u1m_4) + -1.634847819805e-01*V(u1m_5) + 1.830061972141e-01*V(u1m_6)
+ + -2.071774452925e-01*V(u1m_7) + 1.193797886372e-01*V(u1m_8) + 1.082946062088e-01*V(u1m_9) + -1.485439538956e-01*V(u1m_10)
+ + -5.762284994125e-02*V(u1m_11) + 2.465304732323e-02*V(u1m_12) + -3.733760118484e-02*V(u1m_13) + 1.912946999073e-02*V(u1m_14)
+ + 1.109873056412e-01*V(u1m_15) + -1.456275284290e-01*V(u1m_16) + -2.220343053341e-01*V(u1m_17) + 7.713854312897e-02*V(u1m_18)
+ + 5.824449658394e-02*V(u1m_19))
B_u2b_2 u2b_2 0 V = tanh_psi(-3.378880620003e-01 + 1.110349297523e-01*V(u1p_0) + 3.986474871635e-02*V(u1p_1) + 2.204366326332e-01*V(u1p_2)
+ + 1.056722402573e-01*V(u1p_3) + -1.978406906128e-01*V(u1p_4) + -1.634847819805e-01*V(u1p_5) + 1.830061972141e-01*V(u1p_6)
+ + -2.071774452925e-01*V(u1p_7) + 1.193797886372e-01*V(u1p_8) + 1.082946062088e-01*V(u1p_9) + -1.485439538956e-01*V(u1p_10)
+ + -5.762284994125e-02*V(u1p_11) + 2.465304732323e-02*V(u1p_12) + -3.733760118484e-02*V(u1p_13) + 1.912946999073e-02*V(u1p_14)
+ + 1.109873056412e-01*V(u1p_15) + -1.456275284290e-01*V(u1p_16) + -2.220343053341e-01*V(u1p_17) + 7.713854312897e-02*V(u1p_18)
+ + 5.824449658394e-02*V(u1p_19) + 1.407382786274e-01*V(u1m_0) + 2.002112567425e-01*V(u1m_1) + 7.116436958313e-03*V(u1m_2)
+ + 2.026466131210e-01*V(u1m_3) + -8.188287913799e-02*V(u1m_4) + 3.207176923752e-03*V(u1m_5) + -3.131516277790e-02*V(u1m_6)
+ + 1.129356324673e-01*V(u1m_7) + -1.737996488810e-01*V(u1m_8) + 1.128564178944e-01*V(u1m_9) + 8.042323589325e-02*V(u1m_10)
+ + 3.867527842522e-02*V(u1m_11) + -1.359773874283e-01*V(u1m_12) + 1.179875731468e-01*V(u1m_13) + 9.016263484955e-02*V(u1m_14)
+ + -2.096267789602e-01*V(u1m_15) + -1.058997288346e-01*V(u1m_16) + -1.962925493717e-01*V(u1m_17) + -1.598631441593e-01*V(u1m_18)
+ + 7.738000154495e-02*V(u1m_19))
B_u2c_2 u2c_2 0 V = tanh_psi(0.0 + 6.124764680862e-02*(V(u1p_0) + (-1)*V(u1m_0)) + -1.290554106236e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + 9.638306498528e-02*(V(u1p_2) + (-1)*V(u1m_2)) + -1.919362545013e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.335945129395e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 6.839534640312e-02*(V(u1p_5) + (-1)*V(u1m_5)) + 1.334485411644e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + 1.524864733219e-01*(V(u1p_7) + (-1)*V(u1m_7)) + 1.983577013016e-02*(V(u1p_8) + (-1)*V(u1m_8)) + 1.802118420601e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -1.151502430439e-01*(V(u1p_10) + (-1)*V(u1m_10)) + -1.974258273840e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + 1.852292716503e-01*(V(u1p_12) + (-1)*V(u1m_12)) + -1.913675814867e-01*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.564226448536e-01*(V(u1p_14) + (-1)*V(u1m_14)) + -1.391619443893e-02*(V(u1p_15) + (-1)*V(u1m_15))
+ + 4.868423938751e-02*(V(u1p_16) + (-1)*V(u1m_16)) + -2.148323357105e-01*(V(u1p_17) + (-1)*V(u1m_17))
+ + -1.036764308810e-01*(V(u1p_18) + (-1)*V(u1m_18)) + 2.038292586803e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_3 u2a_3 0 V = tanh_psi(9.948115050793e-02 + -1.399420648813e-01*V(u1p_0) + -1.835140883923e-01*V(u1p_1) + 1.384288966656e-01*V(u1p_2)
+ + -2.405913174152e-02*V(u1p_3) + -6.726081669331e-02*V(u1p_4) + -1.608969420195e-01*V(u1p_5) + -4.373027384281e-02*V(u1p_6)
+ + 5.498793721199e-02*V(u1p_7) + 7.528501749039e-02*V(u1p_8) + 4.178142547607e-02*V(u1p_9) + 1.189029514790e-01*V(u1p_10)
+ + -1.862311512232e-01*V(u1p_11) + 3.934293985367e-02*V(u1p_12) + 2.188123464584e-01*V(u1p_13) + 1.203055083752e-01*V(u1p_14)
+ + -4.554453492165e-02*V(u1p_15) + 3.106734156609e-02*V(u1p_16) + 5.294907093048e-02*V(u1p_17) + -2.081075012684e-01*V(u1p_18)
+ + 6.909126043320e-02*V(u1p_19) + -2.837169170380e-02*V(u1m_0) + -1.935914158821e-03*V(u1m_1) + 9.887725114822e-03*V(u1m_2)
+ + -1.430556774139e-01*V(u1m_3) + -1.591846346855e-03*V(u1m_4) + -1.309079974890e-01*V(u1m_5) + -8.249637484550e-02*V(u1m_6)
+ + 9.027755260468e-02*V(u1m_7) + -5.999006330967e-02*V(u1m_8) + -9.401299059391e-02*V(u1m_9) + -7.613837718964e-02*V(u1m_10)
+ + 1.024648249149e-01*V(u1m_11) + 1.112237572670e-02*V(u1m_12) + 6.371417641640e-02*V(u1m_13) + 8.655488491058e-04*V(u1m_14)
+ + -8.227282762527e-02*V(u1m_15) + 3.340703248978e-02*V(u1m_16) + 7.592329382896e-02*V(u1m_17) + 1.803723871708e-01*V(u1m_18)
+ + -1.591103672981e-01*V(u1m_19))
B_u2b_3 u2b_3 0 V = tanh_psi(9.948115050793e-02 + -2.837169170380e-02*V(u1p_0) + -1.935914158821e-03*V(u1p_1) + 9.887725114822e-03*V(u1p_2)
+ + -1.430556774139e-01*V(u1p_3) + -1.591846346855e-03*V(u1p_4) + -1.309079974890e-01*V(u1p_5) + -8.249637484550e-02*V(u1p_6)
+ + 9.027755260468e-02*V(u1p_7) + -5.999006330967e-02*V(u1p_8) + -9.401299059391e-02*V(u1p_9) + -7.613837718964e-02*V(u1p_10)
+ + 1.024648249149e-01*V(u1p_11) + 1.112237572670e-02*V(u1p_12) + 6.371417641640e-02*V(u1p_13) + 8.655488491058e-04*V(u1p_14)
+ + -8.227282762527e-02*V(u1p_15) + 3.340703248978e-02*V(u1p_16) + 7.592329382896e-02*V(u1p_17) + 1.803723871708e-01*V(u1p_18)
+ + -1.591103672981e-01*V(u1p_19) + -1.399420648813e-01*V(u1m_0) + -1.835140883923e-01*V(u1m_1) + 1.384288966656e-01*V(u1m_2)
+ + -2.405913174152e-02*V(u1m_3) + -6.726081669331e-02*V(u1m_4) + -1.608969420195e-01*V(u1m_5) + -4.373027384281e-02*V(u1m_6)
+ + 5.498793721199e-02*V(u1m_7) + 7.528501749039e-02*V(u1m_8) + 4.178142547607e-02*V(u1m_9) + 1.189029514790e-01*V(u1m_10)
+ + -1.862311512232e-01*V(u1m_11) + 3.934293985367e-02*V(u1m_12) + 2.188123464584e-01*V(u1m_13) + 1.203055083752e-01*V(u1m_14)
+ + -4.554453492165e-02*V(u1m_15) + 3.106734156609e-02*V(u1m_16) + 5.294907093048e-02*V(u1m_17) + -2.081075012684e-01*V(u1m_18)
+ + 6.909126043320e-02*V(u1m_19))
B_u2c_3 u2c_3 0 V = tanh_psi(0.0 + -1.145619228482e-01*(V(u1p_0) + (-1)*V(u1m_0)) + -2.073505967855e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + 2.319589257240e-02*(V(u1p_2) + (-1)*V(u1m_2)) + -1.205921173096e-03*(V(u1p_3) + (-1)*V(u1m_3)) + 1.391749978065e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + -1.712366491556e-01*(V(u1p_5) + (-1)*V(u1m_5)) + -5.073994398117e-02*(V(u1p_6) + (-1)*V(u1m_6))
+ + 1.835989952087e-01*(V(u1p_7) + (-1)*V(u1m_7)) + 1.058632731438e-01*(V(u1p_8) + (-1)*V(u1m_8)) + -2.102553844452e-05*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -1.754722297192e-01*(V(u1p_10) + (-1)*V(u1m_10)) + -1.170435920358e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + 3.446415066719e-03*(V(u1p_12) + (-1)*V(u1m_12)) + 1.556347608566e-01*(V(u1p_13) + (-1)*V(u1m_13)) + 2.936908602715e-02*(V(u1p_14)
+ + (-1)*V(u1m_14)) + 2.008709013462e-01*(V(u1p_15) + (-1)*V(u1m_15)) + 2.036512792110e-01*(V(u1p_16) + (-1)*V(u1m_16))
+ + 1.088841855526e-01*(V(u1p_17) + (-1)*V(u1m_17)) + -1.334411799908e-01*(V(u1p_18) + (-1)*V(u1m_18)) + 1.081750392914e-01*(V(u1p_19)
+ + (-1)*V(u1m_19)))
B_u2a_4 u2a_4 0 V = tanh_psi(-2.275057137012e-03 + -1.630178987980e-01*V(u1p_0) + 1.717589795589e-01*V(u1p_1) + 1.233820617199e-01*V(u1p_2)
+ + -2.089801877737e-01*V(u1p_3) + -9.854531288147e-02*V(u1p_4) + -5.742371082306e-03*V(u1p_5) + -1.545462012291e-02*V(u1p_6)
+ + -5.160531401634e-02*V(u1p_7) + 3.682047128677e-02*V(u1p_8) + -1.670405119658e-01*V(u1p_9) + 4.633575677872e-02*V(u1p_10)
+ + 7.774201035500e-02*V(u1p_11) + 8.850145339966e-02*V(u1p_12) + -1.470101177692e-01*V(u1p_13) + 8.060887455940e-03*V(u1p_14)
+ + 5.753171443939e-02*V(u1p_15) + 1.447241306305e-01*V(u1p_16) + 1.569468379021e-01*V(u1p_17) + -1.800000220537e-01*V(u1p_18)
+ + 1.513211429119e-02*V(u1p_19) + -2.082751691341e-02*V(u1m_0) + -2.716046571732e-02*V(u1m_1) + 2.419520914555e-02*V(u1m_2)
+ + 1.471550762653e-01*V(u1m_3) + -6.833124160767e-02*V(u1m_4) + 1.556715667248e-01*V(u1m_5) + -6.452353298664e-02*V(u1m_6)
+ + 8.145469427109e-02*V(u1m_7) + -1.397346854210e-01*V(u1m_8) + -3.765435516834e-02*V(u1m_9) + -5.843126773834e-02*V(u1m_10)
+ + -2.078348696232e-01*V(u1m_11) + -4.642122983932e-02*V(u1m_12) + -1.381921470165e-01*V(u1m_13) + 1.616398394108e-01*V(u1m_14)
+ + 1.852681636810e-01*V(u1m_15) + -5.175872147083e-02*V(u1m_16) + 1.402917206287e-01*V(u1m_17) + -2.846406400204e-02*V(u1m_18)
+ + -1.078324764967e-01*V(u1m_19))
B_u2b_4 u2b_4 0 V = tanh_psi(-2.275057137012e-03 + -2.082751691341e-02*V(u1p_0) + -2.716046571732e-02*V(u1p_1) + 2.419520914555e-02*V(u1p_2)
+ + 1.471550762653e-01*V(u1p_3) + -6.833124160767e-02*V(u1p_4) + 1.556715667248e-01*V(u1p_5) + -6.452353298664e-02*V(u1p_6)
+ + 8.145469427109e-02*V(u1p_7) + -1.397346854210e-01*V(u1p_8) + -3.765435516834e-02*V(u1p_9) + -5.843126773834e-02*V(u1p_10)
+ + -2.078348696232e-01*V(u1p_11) + -4.642122983932e-02*V(u1p_12) + -1.381921470165e-01*V(u1p_13) + 1.616398394108e-01*V(u1p_14)
+ + 1.852681636810e-01*V(u1p_15) + -5.175872147083e-02*V(u1p_16) + 1.402917206287e-01*V(u1p_17) + -2.846406400204e-02*V(u1p_18)
+ + -1.078324764967e-01*V(u1p_19) + -1.630178987980e-01*V(u1m_0) + 1.717589795589e-01*V(u1m_1) + 1.233820617199e-01*V(u1m_2)
+ + -2.089801877737e-01*V(u1m_3) + -9.854531288147e-02*V(u1m_4) + -5.742371082306e-03*V(u1m_5) + -1.545462012291e-02*V(u1m_6)
+ + -5.160531401634e-02*V(u1m_7) + 3.682047128677e-02*V(u1m_8) + -1.670405119658e-01*V(u1m_9) + 4.633575677872e-02*V(u1m_10)
+ + 7.774201035500e-02*V(u1m_11) + 8.850145339966e-02*V(u1m_12) + -1.470101177692e-01*V(u1m_13) + 8.060887455940e-03*V(u1m_14)
+ + 5.753171443939e-02*V(u1m_15) + 1.447241306305e-01*V(u1m_16) + 1.569468379021e-01*V(u1m_17) + -1.800000220537e-01*V(u1m_18)
+ + 1.513211429119e-02*V(u1m_19))
B_u2c_4 u2c_4 0 V = tanh_psi(0.0 + 7.840067148209e-03*(V(u1p_0) + (-1)*V(u1m_0)) + 1.991811394691e-02*(V(u1p_1) + (-1)*V(u1m_1))
+ + 2.198858261108e-01*(V(u1p_2) + (-1)*V(u1m_2)) + -1.613302528858e-01*(V(u1p_3) + (-1)*V(u1m_3)) + -1.917336881161e-02*(V(u1p_4)
+ + (-1)*V(u1m_4)) + -4.183225333691e-02*(V(u1p_5) + (-1)*V(u1m_5)) + -1.597276329994e-02*(V(u1p_6) + (-1)*V(u1m_6))
+ + -1.839578151703e-03*(V(u1p_7) + (-1)*V(u1m_7)) + 6.734719872475e-02*(V(u1p_8) + (-1)*V(u1m_8)) + -1.388624161482e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 2.023020386696e-01*(V(u1p_10) + (-1)*V(u1m_10)) + -2.025324553251e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + -1.633864492178e-01*(V(u1p_12) + (-1)*V(u1m_12)) + 1.756389439106e-01*(V(u1p_13) + (-1)*V(u1m_13)) + 9.457984566689e-02*(V(u1p_14)
+ + (-1)*V(u1m_14)) + 1.013972461224e-01*(V(u1p_15) + (-1)*V(u1m_15)) + -1.337296962738e-01*(V(u1p_16) + (-1)*V(u1m_16))
+ + -2.885347604752e-02*(V(u1p_17) + (-1)*V(u1m_17)) + -1.750712096691e-01*(V(u1p_18) + (-1)*V(u1m_18))
+ + 1.229917407036e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_5 u2a_5 0 V = tanh_psi(8.920190483332e-02 + 1.590909659863e-01*V(u1p_0) + 1.193690001965e-01*V(u1p_1) + -6.945867836475e-02*V(u1p_2)
+ + -1.968015134335e-01*V(u1p_3) + -1.233160495758e-01*V(u1p_4) + 2.699759602547e-02*V(u1p_5) + -2.189186215401e-02*V(u1p_6)
+ + 3.114536404610e-03*V(u1p_7) + 2.095932960510e-01*V(u1p_8) + -1.921945065260e-01*V(u1p_9) + -2.025880813599e-01*V(u1p_10)
+ + -7.435029745102e-02*V(u1p_11) + -1.139027997851e-01*V(u1p_12) + 1.145817935467e-01*V(u1p_13) + 1.895754039288e-01*V(u1p_14)
+ + 5.069914460182e-02*V(u1p_15) + 2.311255037785e-02*V(u1p_16) + -1.218006014824e-01*V(u1p_17) + -4.891987144947e-02*V(u1p_18)
+ + -5.709558725357e-03*V(u1p_19) + -1.616370081902e-01*V(u1m_0) + -1.319043934345e-01*V(u1m_1) + 9.780377149582e-03*V(u1m_2)
+ + -1.079576313496e-01*V(u1m_3) + 7.470050454140e-02*V(u1m_4) + 1.132261753082e-01*V(u1m_5) + 6.370067596436e-02*V(u1m_6)
+ + 5.680900812149e-02*V(u1m_7) + -3.898502886295e-02*V(u1m_8) + -1.183806881309e-01*V(u1m_9) + 4.438728094101e-02*V(u1m_10)
+ + 1.909587681293e-01*V(u1m_11) + -1.333417445421e-01*V(u1m_12) + -1.701995730400e-01*V(u1m_13) + 1.697176694870e-01*V(u1m_14)
+ + -9.729440510273e-02*V(u1m_15) + 1.307555735111e-01*V(u1m_16) + 1.113626956940e-01*V(u1m_17) + -2.162263393402e-01*V(u1m_18)
+ + 1.284810006618e-01*V(u1m_19))
B_u2b_5 u2b_5 0 V = tanh_psi(8.920190483332e-02 + -1.616370081902e-01*V(u1p_0) + -1.319043934345e-01*V(u1p_1) + 9.780377149582e-03*V(u1p_2)
+ + -1.079576313496e-01*V(u1p_3) + 7.470050454140e-02*V(u1p_4) + 1.132261753082e-01*V(u1p_5) + 6.370067596436e-02*V(u1p_6)
+ + 5.680900812149e-02*V(u1p_7) + -3.898502886295e-02*V(u1p_8) + -1.183806881309e-01*V(u1p_9) + 4.438728094101e-02*V(u1p_10)
+ + 1.909587681293e-01*V(u1p_11) + -1.333417445421e-01*V(u1p_12) + -1.701995730400e-01*V(u1p_13) + 1.697176694870e-01*V(u1p_14)
+ + -9.729440510273e-02*V(u1p_15) + 1.307555735111e-01*V(u1p_16) + 1.113626956940e-01*V(u1p_17) + -2.162263393402e-01*V(u1p_18)
+ + 1.284810006618e-01*V(u1p_19) + 1.590909659863e-01*V(u1m_0) + 1.193690001965e-01*V(u1m_1) + -6.945867836475e-02*V(u1m_2)
+ + -1.968015134335e-01*V(u1m_3) + -1.233160495758e-01*V(u1m_4) + 2.699759602547e-02*V(u1m_5) + -2.189186215401e-02*V(u1m_6)
+ + 3.114536404610e-03*V(u1m_7) + 2.095932960510e-01*V(u1m_8) + -1.921945065260e-01*V(u1m_9) + -2.025880813599e-01*V(u1m_10)
+ + -7.435029745102e-02*V(u1m_11) + -1.139027997851e-01*V(u1m_12) + 1.145817935467e-01*V(u1m_13) + 1.895754039288e-01*V(u1m_14)
+ + 5.069914460182e-02*V(u1m_15) + 2.311255037785e-02*V(u1m_16) + -1.218006014824e-01*V(u1m_17) + -4.891987144947e-02*V(u1m_18)
+ + -5.709558725357e-03*V(u1m_19))
B_u2c_5 u2c_5 0 V = tanh_psi(0.0 + 4.828423261642e-04*(V(u1p_0) + (-1)*V(u1m_0)) + -1.799495518208e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + 2.151696383953e-02*(V(u1p_2) + (-1)*V(u1m_2)) + 5.355247855186e-02*(V(u1p_3) + (-1)*V(u1m_3)) + -2.011897563934e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 1.667737960815e-03*(V(u1p_5) + (-1)*V(u1m_5)) + 1.841225624084e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + 1.136304736137e-01*(V(u1p_7) + (-1)*V(u1m_7)) + 6.010705232620e-02*(V(u1p_8) + (-1)*V(u1m_8)) + 2.077549099922e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 1.816636025906e-01*(V(u1p_10) + (-1)*V(u1m_10)) + 9.082794189453e-02*(V(u1p_11) + (-1)*V(u1m_11))
+ + -5.072979629040e-02*(V(u1p_12) + (-1)*V(u1m_12)) + 2.163156569004e-01*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.315108537674e-01*(V(u1p_14) + (-1)*V(u1m_14)) + 1.582274436951e-01*(V(u1p_15) + (-1)*V(u1m_15))
+ + -1.263725012541e-01*(V(u1p_16) + (-1)*V(u1m_16)) + 4.938986897469e-02*(V(u1p_17) + (-1)*V(u1m_17)) + 2.071325182915e-01*(V(u1p_18)
+ + (-1)*V(u1m_18)) + -1.980351209641e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_6 u2a_6 0 V = tanh_psi(-1.041894257069e-01 + -1.661926805973e-01*V(u1p_0) + -5.197022855282e-02*V(u1p_1) + -1.052182689309e-01*V(u1p_2)
+ + 1.889198422432e-01*V(u1p_3) + 4.153260588646e-02*V(u1p_4) + 6.095170974731e-02*V(u1p_5) + 1.381961405277e-01*V(u1p_6)
+ + 2.103078365326e-01*V(u1p_7) + -4.820735752583e-02*V(u1p_8) + 1.871013641357e-01*V(u1p_9) + -2.170673012733e-01*V(u1p_10)
+ + 1.082384884357e-01*V(u1p_11) + 2.674138545990e-02*V(u1p_12) + -1.099959313869e-01*V(u1p_13) + 6.145006418228e-02*V(u1p_14)
+ + 9.870526194572e-02*V(u1p_15) + -5.137257277966e-02*V(u1p_16) + -1.279223859310e-01*V(u1p_17) + 7.450059056282e-03*V(u1p_18)
+ + 1.661272644997e-01*V(u1p_19) + -1.684437692165e-01*V(u1m_0) + 1.968482136726e-01*V(u1m_1) + 1.998093724251e-01*V(u1m_2)
+ + 1.482627987862e-01*V(u1m_3) + 1.235547661781e-01*V(u1m_4) + 1.588805913925e-01*V(u1m_5) + -1.080792844296e-01*V(u1m_6)
+ + -1.901612579823e-01*V(u1m_7) + 1.793685555458e-02*V(u1m_8) + 1.618680357933e-01*V(u1m_9) + -1.166970953345e-01*V(u1m_10)
+ + -5.108679831028e-02*V(u1m_11) + -2.190524786711e-01*V(u1m_12) + 6.643739342690e-02*V(u1m_13) + -1.070348247886e-01*V(u1m_14)
+ + -1.807824075222e-01*V(u1m_15) + -1.195247471333e-02*V(u1m_16) + -1.368078291416e-01*V(u1m_17) + 1.726339161396e-01*V(u1m_18)
+ + -1.218271479011e-01*V(u1m_19))
B_u2b_6 u2b_6 0 V = tanh_psi(-1.041894257069e-01 + -1.684437692165e-01*V(u1p_0) + 1.968482136726e-01*V(u1p_1) + 1.998093724251e-01*V(u1p_2)
+ + 1.482627987862e-01*V(u1p_3) + 1.235547661781e-01*V(u1p_4) + 1.588805913925e-01*V(u1p_5) + -1.080792844296e-01*V(u1p_6)
+ + -1.901612579823e-01*V(u1p_7) + 1.793685555458e-02*V(u1p_8) + 1.618680357933e-01*V(u1p_9) + -1.166970953345e-01*V(u1p_10)
+ + -5.108679831028e-02*V(u1p_11) + -2.190524786711e-01*V(u1p_12) + 6.643739342690e-02*V(u1p_13) + -1.070348247886e-01*V(u1p_14)
+ + -1.807824075222e-01*V(u1p_15) + -1.195247471333e-02*V(u1p_16) + -1.368078291416e-01*V(u1p_17) + 1.726339161396e-01*V(u1p_18)
+ + -1.218271479011e-01*V(u1p_19) + -1.661926805973e-01*V(u1m_0) + -5.197022855282e-02*V(u1m_1) + -1.052182689309e-01*V(u1m_2)
+ + 1.889198422432e-01*V(u1m_3) + 4.153260588646e-02*V(u1m_4) + 6.095170974731e-02*V(u1m_5) + 1.381961405277e-01*V(u1m_6)
+ + 2.103078365326e-01*V(u1m_7) + -4.820735752583e-02*V(u1m_8) + 1.871013641357e-01*V(u1m_9) + -2.170673012733e-01*V(u1m_10)
+ + 1.082384884357e-01*V(u1m_11) + 2.674138545990e-02*V(u1m_12) + -1.099959313869e-01*V(u1m_13) + 6.145006418228e-02*V(u1m_14)
+ + 9.870526194572e-02*V(u1m_15) + -5.137257277966e-02*V(u1m_16) + -1.279223859310e-01*V(u1m_17) + 7.450059056282e-03*V(u1m_18)
+ + 1.661272644997e-01*V(u1m_19))
B_u2c_6 u2c_6 0 V = tanh_psi(0.0 + 1.681973040104e-01*(V(u1p_0) + (-1)*V(u1m_0)) + -1.275362074375e-02*(V(u1p_1) + (-1)*V(u1m_1))
+ + -5.917358398438e-02*(V(u1p_2) + (-1)*V(u1m_2)) + -2.097769677639e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.913412809372e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 1.731294989586e-01*(V(u1p_5) + (-1)*V(u1m_5)) + 1.032012999058e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + 1.876822412014e-01*(V(u1p_7) + (-1)*V(u1m_7)) + -1.914885640144e-01*(V(u1p_8) + (-1)*V(u1m_8)) + 1.433855593204e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -2.008053660393e-02*(V(u1p_10) + (-1)*V(u1m_10)) + 1.653578579426e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + -1.328687071800e-01*(V(u1p_12) + (-1)*V(u1m_12)) + 1.722208857536e-01*(V(u1p_13) + (-1)*V(u1m_13)) + 2.086169421673e-01*(V(u1p_14)
+ + (-1)*V(u1m_14)) + -2.148263305426e-01*(V(u1p_15) + (-1)*V(u1m_15)) + -1.685001403093e-01*(V(u1p_16) + (-1)*V(u1m_16))
+ + 2.217163443565e-01*(V(u1p_17) + (-1)*V(u1m_17)) + -1.079391315579e-01*(V(u1p_18) + (-1)*V(u1m_18))
+ + -1.043182015419e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_7 u2a_7 0 V = tanh_psi(-8.420604467392e-02 + -1.369113326073e-01*V(u1p_0) + 6.994816660881e-02*V(u1p_1) + -7.478228211403e-02*V(u1p_2)
+ + 2.194235920906e-01*V(u1p_3) + -1.034921407700e-02*V(u1p_4) + 2.043696939945e-01*V(u1p_5) + 8.097034692764e-02*V(u1p_6)
+ + -1.893415153027e-01*V(u1p_7) + -2.192481905222e-01*V(u1p_8) + -1.674234867096e-02*V(u1p_9) + 1.038785278797e-01*V(u1p_10)
+ + 1.105797290802e-02*V(u1p_11) + -5.800822377205e-02*V(u1p_12) + -2.613981068134e-02*V(u1p_13) + -5.238375067711e-02*V(u1p_14)
+ + -1.552642881870e-01*V(u1p_15) + -9.332561492920e-02*V(u1p_16) + 1.991002857685e-01*V(u1p_17) + -1.398488283157e-01*V(u1p_18)
+ + -2.389644086361e-02*V(u1p_19) + -9.439563751221e-02*V(u1m_0) + 1.725149452686e-01*V(u1m_1) + 8.424857258797e-02*V(u1m_2)
+ + 1.777112185955e-01*V(u1m_3) + -6.293107569218e-02*V(u1m_4) + -6.081119179726e-03*V(u1m_5) + 1.594874262810e-02*V(u1m_6)
+ + -7.456791400909e-02*V(u1m_7) + 2.660197019577e-02*V(u1m_8) + -1.616796106100e-01*V(u1m_9) + -5.437998473644e-02*V(u1m_10)
+ + -2.082072943449e-01*V(u1m_11) + -1.314023137093e-02*V(u1m_12) + 1.700026988983e-01*V(u1m_13) + -1.162816882133e-01*V(u1m_14)
+ + -8.432553708553e-02*V(u1m_15) + -5.369548499584e-02*V(u1m_16) + -8.524556457996e-02*V(u1m_17) + -3.931324183941e-02*V(u1m_18)
+ + 3.426325321198e-02*V(u1m_19))
B_u2b_7 u2b_7 0 V = tanh_psi(-8.420604467392e-02 + -9.439563751221e-02*V(u1p_0) + 1.725149452686e-01*V(u1p_1) + 8.424857258797e-02*V(u1p_2)
+ + 1.777112185955e-01*V(u1p_3) + -6.293107569218e-02*V(u1p_4) + -6.081119179726e-03*V(u1p_5) + 1.594874262810e-02*V(u1p_6)
+ + -7.456791400909e-02*V(u1p_7) + 2.660197019577e-02*V(u1p_8) + -1.616796106100e-01*V(u1p_9) + -5.437998473644e-02*V(u1p_10)
+ + -2.082072943449e-01*V(u1p_11) + -1.314023137093e-02*V(u1p_12) + 1.700026988983e-01*V(u1p_13) + -1.162816882133e-01*V(u1p_14)
+ + -8.432553708553e-02*V(u1p_15) + -5.369548499584e-02*V(u1p_16) + -8.524556457996e-02*V(u1p_17) + -3.931324183941e-02*V(u1p_18)
+ + 3.426325321198e-02*V(u1p_19) + -1.369113326073e-01*V(u1m_0) + 6.994816660881e-02*V(u1m_1) + -7.478228211403e-02*V(u1m_2)
+ + 2.194235920906e-01*V(u1m_3) + -1.034921407700e-02*V(u1m_4) + 2.043696939945e-01*V(u1m_5) + 8.097034692764e-02*V(u1m_6)
+ + -1.893415153027e-01*V(u1m_7) + -2.192481905222e-01*V(u1m_8) + -1.674234867096e-02*V(u1m_9) + 1.038785278797e-01*V(u1m_10)
+ + 1.105797290802e-02*V(u1m_11) + -5.800822377205e-02*V(u1m_12) + -2.613981068134e-02*V(u1m_13) + -5.238375067711e-02*V(u1m_14)
+ + -1.552642881870e-01*V(u1m_15) + -9.332561492920e-02*V(u1m_16) + 1.991002857685e-01*V(u1m_17) + -1.398488283157e-01*V(u1m_18)
+ + -2.389644086361e-02*V(u1m_19))
B_u2c_7 u2c_7 0 V = tanh_psi(0.0 + -1.405377238989e-01*(V(u1p_0) + (-1)*V(u1m_0)) + -1.466567218304e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + 1.212934851646e-01*(V(u1p_2) + (-1)*V(u1m_2)) + 1.281414330006e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 8.448171615601e-02*(V(u1p_4)
+ + (-1)*V(u1m_4)) + -8.862099051476e-02*(V(u1p_5) + (-1)*V(u1m_5)) + -1.188652962446e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + 1.622685194016e-01*(V(u1p_7) + (-1)*V(u1m_7)) + -2.221408486366e-01*(V(u1p_8) + (-1)*V(u1m_8)) + 7.552310824394e-03*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 9.442189335823e-02*(V(u1p_10) + (-1)*V(u1m_10)) + -7.405182719231e-02*(V(u1p_11) + (-1)*V(u1m_11))
+ + 2.088730931282e-01*(V(u1p_12) + (-1)*V(u1m_12)) + 1.003791391850e-01*(V(u1p_13) + (-1)*V(u1m_13)) + 4.162451624870e-02*(V(u1p_14)
+ + (-1)*V(u1m_14)) + 1.317308843136e-01*(V(u1p_15) + (-1)*V(u1m_15)) + -8.332446217537e-02*(V(u1p_16) + (-1)*V(u1m_16))
+ + -4.173532128334e-03*(V(u1p_17) + (-1)*V(u1m_17)) + 1.073086261749e-01*(V(u1p_18) + (-1)*V(u1m_18)) + 8.399754762650e-03*(V(u1p_19)
+ + (-1)*V(u1m_19)))
B_u2a_8 u2a_8 0 V = tanh_psi(-1.338502019644e-01 + -9.393706917763e-02*V(u1p_0) + 9.605872631073e-02*V(u1p_1) + 1.713530123234e-01*V(u1p_2)
+ + -9.638628363609e-02*V(u1p_3) + -1.946542114019e-01*V(u1p_4) + 6.560009717941e-02*V(u1p_5) + -1.903071999550e-03*V(u1p_6)
+ + -3.326213359833e-02*V(u1p_7) + 2.083002030849e-02*V(u1p_8) + -8.914986252785e-02*V(u1p_9) + -2.217747569084e-01*V(u1p_10)
+ + 1.457785069942e-01*V(u1p_11) + 1.050862371922e-01*V(u1p_12) + 9.140551090240e-03*V(u1p_13) + 2.086980044842e-01*V(u1p_14)
+ + -3.599850833416e-02*V(u1p_15) + -1.372568011284e-01*V(u1p_16) + -2.166361957788e-01*V(u1p_17) + 4.907062649727e-02*V(u1p_18)
+ + 1.513930857182e-01*V(u1p_19) + -1.460992097855e-01*V(u1m_0) + 4.001402854919e-02*V(u1m_1) + 1.277881264687e-01*V(u1m_2)
+ + -3.206586837769e-02*V(u1m_3) + -1.090445518494e-01*V(u1m_4) + 8.840993046761e-03*V(u1m_5) + 1.483240425587e-01*V(u1m_6)
+ + 1.819646060467e-01*V(u1m_7) + -9.246580302715e-02*V(u1m_8) + 6.015974283218e-02*V(u1m_9) + 2.116607725620e-01*V(u1m_10)
+ + -1.729969084263e-01*V(u1m_11) + -1.413109302521e-01*V(u1m_12) + -8.555887639523e-02*V(u1m_13) + -1.053985208273e-01*V(u1m_14)
+ + 6.035700440407e-03*V(u1m_15) + -1.226016357541e-01*V(u1m_16) + -1.764893531799e-03*V(u1m_17) + 1.076755523682e-01*V(u1m_18)
+ + -5.778193473816e-03*V(u1m_19))
B_u2b_8 u2b_8 0 V = tanh_psi(-1.338502019644e-01 + -1.460992097855e-01*V(u1p_0) + 4.001402854919e-02*V(u1p_1) + 1.277881264687e-01*V(u1p_2)
+ + -3.206586837769e-02*V(u1p_3) + -1.090445518494e-01*V(u1p_4) + 8.840993046761e-03*V(u1p_5) + 1.483240425587e-01*V(u1p_6)
+ + 1.819646060467e-01*V(u1p_7) + -9.246580302715e-02*V(u1p_8) + 6.015974283218e-02*V(u1p_9) + 2.116607725620e-01*V(u1p_10)
+ + -1.729969084263e-01*V(u1p_11) + -1.413109302521e-01*V(u1p_12) + -8.555887639523e-02*V(u1p_13) + -1.053985208273e-01*V(u1p_14)
+ + 6.035700440407e-03*V(u1p_15) + -1.226016357541e-01*V(u1p_16) + -1.764893531799e-03*V(u1p_17) + 1.076755523682e-01*V(u1p_18)
+ + -5.778193473816e-03*V(u1p_19) + -9.393706917763e-02*V(u1m_0) + 9.605872631073e-02*V(u1m_1) + 1.713530123234e-01*V(u1m_2)
+ + -9.638628363609e-02*V(u1m_3) + -1.946542114019e-01*V(u1m_4) + 6.560009717941e-02*V(u1m_5) + -1.903071999550e-03*V(u1m_6)
+ + -3.326213359833e-02*V(u1m_7) + 2.083002030849e-02*V(u1m_8) + -8.914986252785e-02*V(u1m_9) + -2.217747569084e-01*V(u1m_10)
+ + 1.457785069942e-01*V(u1m_11) + 1.050862371922e-01*V(u1m_12) + 9.140551090240e-03*V(u1m_13) + 2.086980044842e-01*V(u1m_14)
+ + -3.599850833416e-02*V(u1m_15) + -1.372568011284e-01*V(u1m_16) + -2.166361957788e-01*V(u1m_17) + 4.907062649727e-02*V(u1m_18)
+ + 1.513930857182e-01*V(u1m_19))
B_u2c_8 u2c_8 0 V = tanh_psi(0.0 + -1.708858013153e-01*(V(u1p_0) + (-1)*V(u1m_0)) + 2.765387296677e-02*(V(u1p_1) + (-1)*V(u1m_1))
+ + -1.795759797096e-01*(V(u1p_2) + (-1)*V(u1m_2)) + -1.971129179001e-01*(V(u1p_3) + (-1)*V(u1m_3)) + -9.407795965672e-02*(V(u1p_4)
+ + (-1)*V(u1m_4)) + -1.191918551922e-02*(V(u1p_5) + (-1)*V(u1m_5)) + -9.685859084129e-03*(V(u1p_6) + (-1)*V(u1m_6))
+ + -1.792630851269e-01*(V(u1p_7) + (-1)*V(u1m_7)) + 1.818826794624e-02*(V(u1p_8) + (-1)*V(u1m_8)) + 3.159359097481e-02*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 1.168403029442e-01*(V(u1p_10) + (-1)*V(u1m_10)) + 1.080146133900e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + 7.255417108536e-02*(V(u1p_12) + (-1)*V(u1m_12)) + -5.042447149754e-02*(V(u1p_13) + (-1)*V(u1m_13))
+ + -9.933880716562e-02*(V(u1p_14) + (-1)*V(u1m_14)) + -1.712510883808e-01*(V(u1p_15) + (-1)*V(u1m_15))
+ + 1.158885061741e-01*(V(u1p_16) + (-1)*V(u1m_16)) + 1.345527172089e-01*(V(u1p_17) + (-1)*V(u1m_17)) + 2.047191560268e-01*(V(u1p_18)
+ + (-1)*V(u1m_18)) + 1.643763184547e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_9 u2a_9 0 V = tanh_psi(2.093332260847e-01 + 9.274685382843e-02*V(u1p_0) + -1.027793809772e-01*V(u1p_1) + -2.875140309334e-02*V(u1p_2)
+ + 9.177923202515e-04*V(u1p_3) + -2.201976478100e-01*V(u1p_4) + 1.709846854210e-01*V(u1p_5) + -1.850116997957e-01*V(u1p_6)
+ + 2.940198779106e-02*V(u1p_7) + -2.193342894316e-01*V(u1p_8) + -1.970384120941e-01*V(u1p_9) + -6.207495927811e-03*V(u1p_10)
+ + 1.205378472805e-01*V(u1p_11) + -2.203446626663e-01*V(u1p_12) + -1.481102705002e-01*V(u1p_13) + -9.884951263666e-02*V(u1p_14)
+ + -6.106711924076e-02*V(u1p_15) + -1.296158432961e-01*V(u1p_16) + -1.931240856647e-01*V(u1p_17) + -4.551827907562e-03*V(u1p_18)
+ + 1.540635526180e-01*V(u1p_19) + 1.242372691631e-01*V(u1m_0) + 7.964980602264e-02*V(u1m_1) + 1.066378057003e-01*V(u1m_2)
+ + -1.222652643919e-01*V(u1m_3) + -2.056933939457e-01*V(u1m_4) + 2.082702517509e-02*V(u1m_5) + -9.197413921356e-03*V(u1m_6)
+ + 2.053734362125e-01*V(u1m_7) + -1.637641936541e-01*V(u1m_8) + 1.681575477123e-01*V(u1m_9) + 9.421831369400e-02*V(u1m_10)
+ + -7.327744364738e-02*V(u1m_11) + 1.691852211952e-01*V(u1m_12) + -9.241269528866e-02*V(u1m_13) + 1.442748010159e-01*V(u1m_14)
+ + 2.183824777603e-01*V(u1m_15) + -4.110977053642e-02*V(u1m_16) + 5.987325310707e-02*V(u1m_17) + 1.438866257668e-01*V(u1m_18)
+ + -1.499491631985e-01*V(u1m_19))
B_u2b_9 u2b_9 0 V = tanh_psi(2.093332260847e-01 + 1.242372691631e-01*V(u1p_0) + 7.964980602264e-02*V(u1p_1) + 1.066378057003e-01*V(u1p_2)
+ + -1.222652643919e-01*V(u1p_3) + -2.056933939457e-01*V(u1p_4) + 2.082702517509e-02*V(u1p_5) + -9.197413921356e-03*V(u1p_6)
+ + 2.053734362125e-01*V(u1p_7) + -1.637641936541e-01*V(u1p_8) + 1.681575477123e-01*V(u1p_9) + 9.421831369400e-02*V(u1p_10)
+ + -7.327744364738e-02*V(u1p_11) + 1.691852211952e-01*V(u1p_12) + -9.241269528866e-02*V(u1p_13) + 1.442748010159e-01*V(u1p_14)
+ + 2.183824777603e-01*V(u1p_15) + -4.110977053642e-02*V(u1p_16) + 5.987325310707e-02*V(u1p_17) + 1.438866257668e-01*V(u1p_18)
+ + -1.499491631985e-01*V(u1p_19) + 9.274685382843e-02*V(u1m_0) + -1.027793809772e-01*V(u1m_1) + -2.875140309334e-02*V(u1m_2)
+ + 9.177923202515e-04*V(u1m_3) + -2.201976478100e-01*V(u1m_4) + 1.709846854210e-01*V(u1m_5) + -1.850116997957e-01*V(u1m_6)
+ + 2.940198779106e-02*V(u1m_7) + -2.193342894316e-01*V(u1m_8) + -1.970384120941e-01*V(u1m_9) + -6.207495927811e-03*V(u1m_10)
+ + 1.205378472805e-01*V(u1m_11) + -2.203446626663e-01*V(u1m_12) + -1.481102705002e-01*V(u1m_13) + -9.884951263666e-02*V(u1m_14)
+ + -6.106711924076e-02*V(u1m_15) + -1.296158432961e-01*V(u1m_16) + -1.931240856647e-01*V(u1m_17) + -4.551827907562e-03*V(u1m_18)
+ + 1.540635526180e-01*V(u1m_19))
B_u2c_9 u2c_9 0 V = tanh_psi(0.0 + 1.108879148960e-01*(V(u1p_0) + (-1)*V(u1m_0)) + -1.939167976379e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + -3.649516403675e-02*(V(u1p_2) + (-1)*V(u1m_2)) + 1.319243013859e-01*(V(u1p_3) + (-1)*V(u1m_3)) + -7.847219705582e-02*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 1.608988642693e-02*(V(u1p_5) + (-1)*V(u1m_5)) + 1.960699558258e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + -1.625729352236e-01*(V(u1p_7) + (-1)*V(u1m_7)) + -1.492415964603e-01*(V(u1p_8) + (-1)*V(u1m_8)) + -5.271206796169e-02*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 2.804455161095e-02*(V(u1p_10) + (-1)*V(u1m_10)) + -6.093406677246e-02*(V(u1p_11) + (-1)*V(u1m_11))
+ + -6.140755116940e-02*(V(u1p_12) + (-1)*V(u1m_12)) + -4.777103662491e-02*(V(u1p_13) + (-1)*V(u1m_13))
+ + 1.749470829964e-02*(V(u1p_14) + (-1)*V(u1m_14)) + 4.590117931366e-02*(V(u1p_15) + (-1)*V(u1m_15)) + 1.385400593281e-01*(V(u1p_16)
+ + (-1)*V(u1m_16)) + -4.528282582760e-02*(V(u1p_17) + (-1)*V(u1m_17)) + 4.410028457642e-02*(V(u1p_18) + (-1)*V(u1m_18))
+ + 1.053055524826e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_10 u2a_10 0 V = tanh_psi(7.425931096077e-02 + -1.563691198826e-01*V(u1p_0) + -1.185403540730e-01*V(u1p_1) + -1.769348978996e-02*V(u1p_2)
+ + -5.121858417988e-02*V(u1p_3) + -1.832500100136e-03*V(u1p_4) + 2.072350084782e-01*V(u1p_5) + 9.344816207886e-04*V(u1p_6)
+ + -2.221954911947e-01*V(u1p_7) + -2.342021465302e-02*V(u1p_8) + 2.198776602745e-01*V(u1p_9) + -4.846736788750e-02*V(u1p_10)
+ + 9.082478284836e-02*V(u1p_11) + 1.390324831009e-01*V(u1p_12) + -2.090690881014e-01*V(u1p_13) + 1.753732264042e-01*V(u1p_14)
+ + -6.522084772587e-02*V(u1p_15) + -5.698801577091e-02*V(u1p_16) + 1.303561925888e-01*V(u1p_17) + 2.058980464935e-01*V(u1p_18)
+ + -2.142037004232e-01*V(u1p_19) + -8.422231674194e-02*V(u1m_0) + -2.051230072975e-01*V(u1m_1) + 1.654741168022e-02*V(u1m_2)
+ + 1.572307050228e-01*V(u1m_3) + 1.414517462254e-01*V(u1m_4) + -7.302783429623e-02*V(u1m_5) + -4.428951442242e-02*V(u1m_6)
+ + -1.226614266634e-01*V(u1m_7) + 1.552324593067e-01*V(u1m_8) + 2.032562196255e-01*V(u1m_9) + -4.793414473534e-02*V(u1m_10)
+ + 1.597528159618e-01*V(u1m_11) + 1.289993524551e-01*V(u1m_12) + 1.409406960011e-01*V(u1m_13) + -8.167307078838e-02*V(u1m_14)
+ + -1.992411911488e-02*V(u1m_15) + -1.371150016785e-01*V(u1m_16) + 2.197290062904e-01*V(u1m_17) + 3.843051195145e-02*V(u1m_18)
+ + -5.613605678082e-02*V(u1m_19))
B_u2b_10 u2b_10 0 V = tanh_psi(7.425931096077e-02 + -8.422231674194e-02*V(u1p_0) + -2.051230072975e-01*V(u1p_1) + 1.654741168022e-02*V(u1p_2)
+ + 1.572307050228e-01*V(u1p_3) + 1.414517462254e-01*V(u1p_4) + -7.302783429623e-02*V(u1p_5) + -4.428951442242e-02*V(u1p_6)
+ + -1.226614266634e-01*V(u1p_7) + 1.552324593067e-01*V(u1p_8) + 2.032562196255e-01*V(u1p_9) + -4.793414473534e-02*V(u1p_10)
+ + 1.597528159618e-01*V(u1p_11) + 1.289993524551e-01*V(u1p_12) + 1.409406960011e-01*V(u1p_13) + -8.167307078838e-02*V(u1p_14)
+ + -1.992411911488e-02*V(u1p_15) + -1.371150016785e-01*V(u1p_16) + 2.197290062904e-01*V(u1p_17) + 3.843051195145e-02*V(u1p_18)
+ + -5.613605678082e-02*V(u1p_19) + -1.563691198826e-01*V(u1m_0) + -1.185403540730e-01*V(u1m_1) + -1.769348978996e-02*V(u1m_2)
+ + -5.121858417988e-02*V(u1m_3) + -1.832500100136e-03*V(u1m_4) + 2.072350084782e-01*V(u1m_5) + 9.344816207886e-04*V(u1m_6)
+ + -2.221954911947e-01*V(u1m_7) + -2.342021465302e-02*V(u1m_8) + 2.198776602745e-01*V(u1m_9) + -4.846736788750e-02*V(u1m_10)
+ + 9.082478284836e-02*V(u1m_11) + 1.390324831009e-01*V(u1m_12) + -2.090690881014e-01*V(u1m_13) + 1.753732264042e-01*V(u1m_14)
+ + -6.522084772587e-02*V(u1m_15) + -5.698801577091e-02*V(u1m_16) + 1.303561925888e-01*V(u1m_17) + 2.058980464935e-01*V(u1m_18)
+ + -2.142037004232e-01*V(u1m_19))
B_u2c_10 u2c_10 0 V = tanh_psi(0.0 + -6.296485662460e-04*(V(u1p_0) + (-1)*V(u1m_0)) + 1.206092238426e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + -2.217453271151e-01*(V(u1p_2) + (-1)*V(u1m_2)) + -1.409113556147e-01*(V(u1p_3) + (-1)*V(u1m_3)) + -1.631464064121e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + -7.720187306404e-03*(V(u1p_5) + (-1)*V(u1m_5)) + 8.337834477425e-02*(V(u1p_6) + (-1)*V(u1m_6))
+ + 6.032705307007e-03*(V(u1p_7) + (-1)*V(u1m_7)) + -1.797525137663e-01*(V(u1p_8) + (-1)*V(u1m_8)) + 1.934753060341e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 7.847800850868e-03*(V(u1p_10) + (-1)*V(u1m_10)) + 1.684336364269e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + 1.725550293922e-01*(V(u1p_12) + (-1)*V(u1m_12)) + -5.464060604572e-02*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.627555787563e-01*(V(u1p_14) + (-1)*V(u1m_14)) + 9.885969758034e-02*(V(u1p_15) + (-1)*V(u1m_15))
+ + -1.125088185072e-01*(V(u1p_16) + (-1)*V(u1m_16)) + -1.558677554131e-01*(V(u1p_17) + (-1)*V(u1m_17))
+ + -8.565513789654e-02*(V(u1p_18) + (-1)*V(u1m_18)) + -1.266588419676e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_11 u2a_11 0 V = tanh_psi(-4.129375517368e-02 + -3.809884190559e-03*V(u1p_0) + 9.487569332123e-02*V(u1p_1) + -1.814135611057e-01*V(u1p_2)
+ + 1.038120985031e-01*V(u1p_3) + 1.677136719227e-01*V(u1p_4) + -2.137550264597e-01*V(u1p_5) + -2.195223420858e-01*V(u1p_6)
+ + 1.716342270374e-01*V(u1p_7) + -1.908286213875e-01*V(u1p_8) + 6.433227658272e-02*V(u1p_9) + -2.033655345440e-01*V(u1p_10)
+ + 1.553535163403e-01*V(u1p_11) + 6.299689412117e-03*V(u1p_12) + -1.349435150623e-01*V(u1p_13) + 1.810340881348e-01*V(u1p_14)
+ + 7.635250687599e-02*V(u1p_15) + 2.096390426159e-01*V(u1p_16) + 1.686590611935e-01*V(u1p_17) + -1.633361726999e-01*V(u1p_18)
+ + -7.751454412937e-02*V(u1p_19) + 6.451240181923e-02*V(u1m_0) + 5.933803319931e-02*V(u1m_1) + -1.767255961895e-01*V(u1m_2)
+ + 1.250684261322e-01*V(u1m_3) + 5.695092678070e-02*V(u1m_4) + -6.286169588566e-02*V(u1m_5) + -1.409557461739e-01*V(u1m_6)
+ + 1.428359746933e-01*V(u1m_7) + -4.001569747925e-02*V(u1m_8) + 2.102590203285e-01*V(u1m_9) + 2.294023334980e-02*V(u1m_10)
+ + 5.804833769798e-02*V(u1m_11) + -6.100504100323e-02*V(u1m_12) + -7.988810539246e-02*V(u1m_13) + 2.010168135166e-01*V(u1m_14)
+ + 1.332529187202e-01*V(u1m_15) + -3.992544114590e-02*V(u1m_16) + -1.929076313972e-01*V(u1m_17) + 1.296983361244e-01*V(u1m_18)
+ + 3.632083535194e-02*V(u1m_19))
B_u2b_11 u2b_11 0 V = tanh_psi(-4.129375517368e-02 + 6.451240181923e-02*V(u1p_0) + 5.933803319931e-02*V(u1p_1) + -1.767255961895e-01*V(u1p_2)
+ + 1.250684261322e-01*V(u1p_3) + 5.695092678070e-02*V(u1p_4) + -6.286169588566e-02*V(u1p_5) + -1.409557461739e-01*V(u1p_6)
+ + 1.428359746933e-01*V(u1p_7) + -4.001569747925e-02*V(u1p_8) + 2.102590203285e-01*V(u1p_9) + 2.294023334980e-02*V(u1p_10)
+ + 5.804833769798e-02*V(u1p_11) + -6.100504100323e-02*V(u1p_12) + -7.988810539246e-02*V(u1p_13) + 2.010168135166e-01*V(u1p_14)
+ + 1.332529187202e-01*V(u1p_15) + -3.992544114590e-02*V(u1p_16) + -1.929076313972e-01*V(u1p_17) + 1.296983361244e-01*V(u1p_18)
+ + 3.632083535194e-02*V(u1p_19) + -3.809884190559e-03*V(u1m_0) + 9.487569332123e-02*V(u1m_1) + -1.814135611057e-01*V(u1m_2)
+ + 1.038120985031e-01*V(u1m_3) + 1.677136719227e-01*V(u1m_4) + -2.137550264597e-01*V(u1m_5) + -2.195223420858e-01*V(u1m_6)
+ + 1.716342270374e-01*V(u1m_7) + -1.908286213875e-01*V(u1m_8) + 6.433227658272e-02*V(u1m_9) + -2.033655345440e-01*V(u1m_10)
+ + 1.553535163403e-01*V(u1m_11) + 6.299689412117e-03*V(u1m_12) + -1.349435150623e-01*V(u1m_13) + 1.810340881348e-01*V(u1m_14)
+ + 7.635250687599e-02*V(u1m_15) + 2.096390426159e-01*V(u1m_16) + 1.686590611935e-01*V(u1m_17) + -1.633361726999e-01*V(u1m_18)
+ + -7.751454412937e-02*V(u1m_19))
B_u2c_11 u2c_11 0 V = tanh_psi(0.0 + -1.016375422478e-02*(V(u1p_0) + (-1)*V(u1m_0)) + 1.959737837315e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + 7.596871256828e-02*(V(u1p_2) + (-1)*V(u1m_2)) + 8.358317613602e-02*(V(u1p_3) + (-1)*V(u1m_3)) + -5.300389230251e-02*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 1.444790065289e-01*(V(u1p_5) + (-1)*V(u1m_5)) + 1.741924285889e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + 3.657114505768e-02*(V(u1p_7) + (-1)*V(u1m_7)) + -1.334526538849e-01*(V(u1p_8) + (-1)*V(u1m_8)) + 1.979252398014e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -1.755087971687e-01*(V(u1p_10) + (-1)*V(u1m_10)) + -1.525730490685e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + -4.398214817047e-02*(V(u1p_12) + (-1)*V(u1m_12)) + -1.162375956774e-01*(V(u1p_13) + (-1)*V(u1m_13))
+ + 1.990455389023e-02*(V(u1p_14) + (-1)*V(u1m_14)) + -2.120501846075e-01*(V(u1p_15) + (-1)*V(u1m_15))
+ + -1.907728016376e-01*(V(u1p_16) + (-1)*V(u1m_16)) + -1.414305269718e-01*(V(u1p_17) + (-1)*V(u1m_17))
+ + 1.458243131638e-01*(V(u1p_18) + (-1)*V(u1m_18)) + -1.253883391619e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_12 u2a_12 0 V = tanh_psi(-1.042537540197e-01 + -4.628111422062e-02*V(u1p_0) + 6.077778339386e-02*V(u1p_1) + 5.583372712135e-02*V(u1p_2)
+ + -1.033079698682e-01*V(u1p_3) + 1.225022673607e-01*V(u1p_4) + 1.201322674751e-01*V(u1p_5) + -8.291639387608e-02*V(u1p_6)
+ + -1.014476194978e-01*V(u1p_7) + 2.094651162624e-01*V(u1p_8) + 1.224400103092e-01*V(u1p_9) + 2.227678894997e-01*V(u1p_10)
+ + 1.861645877361e-01*V(u1p_11) + 6.102880835533e-02*V(u1p_12) + -1.699773967266e-02*V(u1p_13) + -2.092955261469e-01*V(u1p_14)
+ + -5.636863410473e-02*V(u1p_15) + 1.405702531338e-01*V(u1p_16) + 1.121822595596e-01*V(u1p_17) + 4.148602485657e-02*V(u1p_18)
+ + -1.007677838206e-01*V(u1p_19) + -9.814614057541e-02*V(u1m_0) + 2.101570367813e-01*V(u1m_1) + 1.942116022110e-01*V(u1m_2)
+ + -1.559568047523e-01*V(u1m_3) + 9.257844090462e-02*V(u1m_4) + -4.467882215977e-02*V(u1m_5) + -1.785041689873e-01*V(u1m_6)
+ + -1.138029471040e-01*V(u1m_7) + 2.127906680107e-01*V(u1m_8) + 1.297031342983e-02*V(u1m_9) + 1.534643769264e-01*V(u1m_10)
+ + -1.173912733793e-01*V(u1m_11) + -1.556070297956e-01*V(u1m_12) + 4.814440011978e-02*V(u1m_13) + -3.376044332981e-02*V(u1m_14)
+ + 4.836738109589e-02*V(u1m_15) + -1.145347058773e-01*V(u1m_16) + 1.620129346848e-01*V(u1m_17) + 9.361526370049e-02*V(u1m_18)
+ + -3.119941055775e-02*V(u1m_19))
B_u2b_12 u2b_12 0 V = tanh_psi(-1.042537540197e-01 + -9.814614057541e-02*V(u1p_0) + 2.101570367813e-01*V(u1p_1) + 1.942116022110e-01*V(u1p_2)
+ + -1.559568047523e-01*V(u1p_3) + 9.257844090462e-02*V(u1p_4) + -4.467882215977e-02*V(u1p_5) + -1.785041689873e-01*V(u1p_6)
+ + -1.138029471040e-01*V(u1p_7) + 2.127906680107e-01*V(u1p_8) + 1.297031342983e-02*V(u1p_9) + 1.534643769264e-01*V(u1p_10)
+ + -1.173912733793e-01*V(u1p_11) + -1.556070297956e-01*V(u1p_12) + 4.814440011978e-02*V(u1p_13) + -3.376044332981e-02*V(u1p_14)
+ + 4.836738109589e-02*V(u1p_15) + -1.145347058773e-01*V(u1p_16) + 1.620129346848e-01*V(u1p_17) + 9.361526370049e-02*V(u1p_18)
+ + -3.119941055775e-02*V(u1p_19) + -4.628111422062e-02*V(u1m_0) + 6.077778339386e-02*V(u1m_1) + 5.583372712135e-02*V(u1m_2)
+ + -1.033079698682e-01*V(u1m_3) + 1.225022673607e-01*V(u1m_4) + 1.201322674751e-01*V(u1m_5) + -8.291639387608e-02*V(u1m_6)
+ + -1.014476194978e-01*V(u1m_7) + 2.094651162624e-01*V(u1m_8) + 1.224400103092e-01*V(u1m_9) + 2.227678894997e-01*V(u1m_10)
+ + 1.861645877361e-01*V(u1m_11) + 6.102880835533e-02*V(u1m_12) + -1.699773967266e-02*V(u1m_13) + -2.092955261469e-01*V(u1m_14)
+ + -5.636863410473e-02*V(u1m_15) + 1.405702531338e-01*V(u1m_16) + 1.121822595596e-01*V(u1m_17) + 4.148602485657e-02*V(u1m_18)
+ + -1.007677838206e-01*V(u1m_19))
B_u2c_12 u2c_12 0 V = tanh_psi(0.0 + -8.268725872040e-02*(V(u1p_0) + (-1)*V(u1m_0)) + -7.147713005543e-02*(V(u1p_1) + (-1)*V(u1m_1))
+ + 1.111198961735e-01*(V(u1p_2) + (-1)*V(u1m_2)) + 1.460359096527e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.174933314323e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 1.552881002426e-01*(V(u1p_5) + (-1)*V(u1m_5)) + 1.558786928654e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + -2.665907144547e-02*(V(u1p_7) + (-1)*V(u1m_7)) + 2.122578024864e-01*(V(u1p_8) + (-1)*V(u1m_8)) + 1.301470100880e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 1.580953001976e-01*(V(u1p_10) + (-1)*V(u1m_10)) + -2.675679326057e-02*(V(u1p_11) + (-1)*V(u1m_11))
+ + 1.447456777096e-01*(V(u1p_12) + (-1)*V(u1m_12)) + 1.362002789974e-01*(V(u1p_13) + (-1)*V(u1m_13)) + 3.053969144821e-02*(V(u1p_14)
+ + (-1)*V(u1m_14)) + -1.791985034943e-01*(V(u1p_15) + (-1)*V(u1m_15)) + -4.014989733696e-02*(V(u1p_16) + (-1)*V(u1m_16))
+ + 2.981168031693e-02*(V(u1p_17) + (-1)*V(u1m_17)) + -7.232336699963e-02*(V(u1p_18) + (-1)*V(u1m_18))
+ + -6.955876946449e-02*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_13 u2a_13 0 V = tanh_psi(1.942885816097e-01 + 1.256399452686e-01*V(u1p_0) + -1.610043346882e-01*V(u1p_1) + 1.953668594360e-01*V(u1p_2)
+ + -2.080487459898e-01*V(u1p_3) + 3.531408309937e-02*V(u1p_4) + 4.849219322205e-02*V(u1p_5) + -3.523668646812e-02*V(u1p_6)
+ + -7.831713557243e-02*V(u1p_7) + 1.200896501541e-02*V(u1p_8) + 1.408006548882e-01*V(u1p_9) + -1.826577484608e-01*V(u1p_10)
+ + -2.679926156998e-02*V(u1p_11) + 3.493583202362e-02*V(u1p_12) + -1.922760903835e-01*V(u1p_13) + 7.738769054413e-02*V(u1p_14)
+ + -1.979934126139e-01*V(u1p_15) + 1.637312769890e-02*V(u1p_16) + -2.061192095280e-01*V(u1p_17) + -1.186795532703e-01*V(u1p_18)
+ + -1.963968575001e-02*V(u1p_19) + 6.981572508812e-02*V(u1m_0) + -4.695077240467e-02*V(u1m_1) + 1.526216566563e-01*V(u1m_2)
+ + 1.698608398438e-01*V(u1m_3) + -1.918467730284e-01*V(u1m_4) + 1.611513495445e-01*V(u1m_5) + 1.496409773827e-01*V(u1m_6)
+ + 1.865222156048e-01*V(u1m_7) + 3.644213080406e-02*V(u1m_8) + -1.999330073595e-01*V(u1m_9) + -8.951108157635e-02*V(u1m_10)
+ + 1.931017041206e-01*V(u1m_11) + 4.409492015839e-02*V(u1m_12) + -1.036817356944e-01*V(u1m_13) + -2.164832502604e-01*V(u1m_14)
+ + -1.248982697725e-01*V(u1m_15) + 1.976331472397e-01*V(u1m_16) + 1.922486722469e-02*V(u1m_17) + 1.304375231266e-01*V(u1m_18)
+ + 4.348769783974e-03*V(u1m_19))
B_u2b_13 u2b_13 0 V = tanh_psi(1.942885816097e-01 + 6.981572508812e-02*V(u1p_0) + -4.695077240467e-02*V(u1p_1) + 1.526216566563e-01*V(u1p_2)
+ + 1.698608398438e-01*V(u1p_3) + -1.918467730284e-01*V(u1p_4) + 1.611513495445e-01*V(u1p_5) + 1.496409773827e-01*V(u1p_6)
+ + 1.865222156048e-01*V(u1p_7) + 3.644213080406e-02*V(u1p_8) + -1.999330073595e-01*V(u1p_9) + -8.951108157635e-02*V(u1p_10)
+ + 1.931017041206e-01*V(u1p_11) + 4.409492015839e-02*V(u1p_12) + -1.036817356944e-01*V(u1p_13) + -2.164832502604e-01*V(u1p_14)
+ + -1.248982697725e-01*V(u1p_15) + 1.976331472397e-01*V(u1p_16) + 1.922486722469e-02*V(u1p_17) + 1.304375231266e-01*V(u1p_18)
+ + 4.348769783974e-03*V(u1p_19) + 1.256399452686e-01*V(u1m_0) + -1.610043346882e-01*V(u1m_1) + 1.953668594360e-01*V(u1m_2)
+ + -2.080487459898e-01*V(u1m_3) + 3.531408309937e-02*V(u1m_4) + 4.849219322205e-02*V(u1m_5) + -3.523668646812e-02*V(u1m_6)
+ + -7.831713557243e-02*V(u1m_7) + 1.200896501541e-02*V(u1m_8) + 1.408006548882e-01*V(u1m_9) + -1.826577484608e-01*V(u1m_10)
+ + -2.679926156998e-02*V(u1m_11) + 3.493583202362e-02*V(u1m_12) + -1.922760903835e-01*V(u1m_13) + 7.738769054413e-02*V(u1m_14)
+ + -1.979934126139e-01*V(u1m_15) + 1.637312769890e-02*V(u1m_16) + -2.061192095280e-01*V(u1m_17) + -1.186795532703e-01*V(u1m_18)
+ + -1.963968575001e-02*V(u1m_19))
B_u2c_13 u2c_13 0 V = tanh_psi(0.0 + 2.332800626755e-02*(V(u1p_0) + (-1)*V(u1m_0)) + -6.110289692879e-02*(V(u1p_1) + (-1)*V(u1m_1))
+ + -2.213527560234e-01*(V(u1p_2) + (-1)*V(u1m_2)) + 1.712850630283e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.617998182774e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 2.032017707825e-01*(V(u1p_5) + (-1)*V(u1m_5)) + -9.739907085896e-02*(V(u1p_6) + (-1)*V(u1m_6))
+ + 6.207033991814e-03*(V(u1p_7) + (-1)*V(u1m_7)) + 3.486269712448e-02*(V(u1p_8) + (-1)*V(u1m_8)) + 1.953949332237e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 5.689403414726e-02*(V(u1p_10) + (-1)*V(u1m_10)) + -1.002786457539e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + -1.653431057930e-01*(V(u1p_12) + (-1)*V(u1m_12)) + -1.345115602016e-01*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.482025980949e-01*(V(u1p_14) + (-1)*V(u1m_14)) + 8.365416526794e-02*(V(u1p_15) + (-1)*V(u1m_15))
+ + -8.662909269333e-03*(V(u1p_16) + (-1)*V(u1m_16)) + -6.799381971359e-02*(V(u1p_17) + (-1)*V(u1m_17))
+ + -2.181541025639e-01*(V(u1p_18) + (-1)*V(u1m_18)) + 2.089866995811e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_14 u2a_14 0 V = tanh_psi(-1.452559232712e-02 + -9.819880127907e-03*V(u1p_0) + -8.538451790810e-02*V(u1p_1) + -1.129880174994e-01*V(u1p_2)
+ + 1.538450717926e-01*V(u1p_3) + 2.140130102634e-01*V(u1p_4) + -1.646596491337e-01*V(u1p_5) + 1.326317489147e-01*V(u1p_6)
+ + -1.891017705202e-01*V(u1p_7) + 1.146672368050e-01*V(u1p_8) + -2.634315192699e-02*V(u1p_9) + -3.426584601402e-02*V(u1p_10)
+ + -1.434044241905e-01*V(u1p_11) + 6.613877415657e-02*V(u1p_12) + -9.026065468788e-03*V(u1p_13) + 1.703140139580e-01*V(u1p_14)
+ + 2.153912186623e-01*V(u1p_15) + 2.012176811695e-01*V(u1p_16) + -3.256580233574e-02*V(u1p_17) + 1.847726106644e-01*V(u1p_18)
+ + 1.302264630795e-01*V(u1p_19) + 9.694629907608e-02*V(u1m_0) + -2.628993988037e-02*V(u1m_1) + -1.962708234787e-01*V(u1m_2)
+ + 4.905477166176e-03*V(u1m_3) + 6.614986062050e-02*V(u1m_4) + -9.178441762924e-02*V(u1m_5) + 1.709842383862e-01*V(u1m_6)
+ + 1.873828172684e-01*V(u1m_7) + -1.256905496120e-02*V(u1m_8) + 1.347700059414e-01*V(u1m_9) + 1.451078653336e-01*V(u1m_10)
+ + -7.833613455296e-02*V(u1m_11) + 1.379664242268e-02*V(u1m_12) + -1.182852610946e-01*V(u1m_13) + 2.212926745415e-03*V(u1m_14)
+ + -1.846394240856e-01*V(u1m_15) + -4.302407801151e-02*V(u1m_16) + -1.403702646494e-01*V(u1m_17) + -1.788139939308e-01*V(u1m_18)
+ + -5.380688607693e-02*V(u1m_19))
B_u2b_14 u2b_14 0 V = tanh_psi(-1.452559232712e-02 + 9.694629907608e-02*V(u1p_0) + -2.628993988037e-02*V(u1p_1) + -1.962708234787e-01*V(u1p_2)
+ + 4.905477166176e-03*V(u1p_3) + 6.614986062050e-02*V(u1p_4) + -9.178441762924e-02*V(u1p_5) + 1.709842383862e-01*V(u1p_6)
+ + 1.873828172684e-01*V(u1p_7) + -1.256905496120e-02*V(u1p_8) + 1.347700059414e-01*V(u1p_9) + 1.451078653336e-01*V(u1p_10)
+ + -7.833613455296e-02*V(u1p_11) + 1.379664242268e-02*V(u1p_12) + -1.182852610946e-01*V(u1p_13) + 2.212926745415e-03*V(u1p_14)
+ + -1.846394240856e-01*V(u1p_15) + -4.302407801151e-02*V(u1p_16) + -1.403702646494e-01*V(u1p_17) + -1.788139939308e-01*V(u1p_18)
+ + -5.380688607693e-02*V(u1p_19) + -9.819880127907e-03*V(u1m_0) + -8.538451790810e-02*V(u1m_1) + -1.129880174994e-01*V(u1m_2)
+ + 1.538450717926e-01*V(u1m_3) + 2.140130102634e-01*V(u1m_4) + -1.646596491337e-01*V(u1m_5) + 1.326317489147e-01*V(u1m_6)
+ + -1.891017705202e-01*V(u1m_7) + 1.146672368050e-01*V(u1m_8) + -2.634315192699e-02*V(u1m_9) + -3.426584601402e-02*V(u1m_10)
+ + -1.434044241905e-01*V(u1m_11) + 6.613877415657e-02*V(u1m_12) + -9.026065468788e-03*V(u1m_13) + 1.703140139580e-01*V(u1m_14)
+ + 2.153912186623e-01*V(u1m_15) + 2.012176811695e-01*V(u1m_16) + -3.256580233574e-02*V(u1m_17) + 1.847726106644e-01*V(u1m_18)
+ + 1.302264630795e-01*V(u1m_19))
B_u2c_14 u2c_14 0 V = tanh_psi(0.0 + 1.080798506737e-01*(V(u1p_0) + (-1)*V(u1m_0)) + 1.323521435261e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + 1.477892696857e-01*(V(u1p_2) + (-1)*V(u1m_2)) + -2.143488675356e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.461012959480e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 8.234003186226e-02*(V(u1p_5) + (-1)*V(u1m_5)) + 8.094528317451e-02*(V(u1p_6) + (-1)*V(u1m_6))
+ + -2.063126116991e-01*(V(u1p_7) + (-1)*V(u1m_7)) + 1.503062248230e-02*(V(u1p_8) + (-1)*V(u1m_8)) + -1.557357013226e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 9.128198027611e-02*(V(u1p_10) + (-1)*V(u1m_10)) + -1.605147719383e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + -1.562834680080e-01*(V(u1p_12) + (-1)*V(u1m_12)) + -1.956724673510e-01*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.686694622040e-01*(V(u1p_14) + (-1)*V(u1m_14)) + -5.163210630417e-02*(V(u1p_15) + (-1)*V(u1m_15))
+ + -1.581549346447e-01*(V(u1p_16) + (-1)*V(u1m_16)) + 1.347814500332e-01*(V(u1p_17) + (-1)*V(u1m_17)) + 2.443161606789e-02*(V(u1p_18)
+ + (-1)*V(u1m_18)) + -1.031745001674e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_15 u2a_15 0 V = tanh_psi(1.740372180939e-01 + 6.992545723915e-02*V(u1p_0) + -4.322490096092e-02*V(u1p_1) + 1.052170991898e-03*V(u1p_2)
+ + -1.664206534624e-01*V(u1p_3) + -4.050457477570e-02*V(u1p_4) + 1.649064421654e-01*V(u1p_5) + -1.753352582455e-02*V(u1p_6)
+ + 1.747005283833e-01*V(u1p_7) + 1.718393862247e-01*V(u1p_8) + 1.166446208954e-01*V(u1p_9) + -3.587155044079e-02*V(u1p_10)
+ + 1.965202689171e-01*V(u1p_11) + 1.127580404282e-01*V(u1p_12) + -2.177745997906e-01*V(u1p_13) + -2.144685536623e-01*V(u1p_14)
+ + -1.371018588543e-01*V(u1p_15) + -1.702023148537e-01*V(u1p_16) + -1.338601708412e-01*V(u1p_17) + 9.209856390953e-02*V(u1p_18)
+ + -1.849099546671e-01*V(u1p_19) + 2.184267640114e-01*V(u1m_0) + 2.223142385483e-01*V(u1m_1) + -1.441995650530e-01*V(u1m_2)
+ + 1.702958643436e-01*V(u1m_3) + 1.710635423660e-02*V(u1m_4) + 1.303254067898e-01*V(u1m_5) + -2.017352283001e-01*V(u1m_6)
+ + 8.896613121033e-02*V(u1m_7) + 1.877025067806e-01*V(u1m_8) + -5.465331673622e-02*V(u1m_9) + -1.301475465298e-01*V(u1m_10)
+ + 1.321718692780e-01*V(u1m_11) + 2.209012508392e-01*V(u1m_12) + 1.083862483501e-01*V(u1m_13) + 1.289784610271e-01*V(u1m_14)
+ + 1.599046289921e-01*V(u1m_15) + 1.521005928516e-01*V(u1m_16) + -4.721339046955e-02*V(u1m_17) + 5.895599722862e-02*V(u1m_18)
+ + 8.082774281502e-02*V(u1m_19))
B_u2b_15 u2b_15 0 V = tanh_psi(1.740372180939e-01 + 2.184267640114e-01*V(u1p_0) + 2.223142385483e-01*V(u1p_1) + -1.441995650530e-01*V(u1p_2)
+ + 1.702958643436e-01*V(u1p_3) + 1.710635423660e-02*V(u1p_4) + 1.303254067898e-01*V(u1p_5) + -2.017352283001e-01*V(u1p_6)
+ + 8.896613121033e-02*V(u1p_7) + 1.877025067806e-01*V(u1p_8) + -5.465331673622e-02*V(u1p_9) + -1.301475465298e-01*V(u1p_10)
+ + 1.321718692780e-01*V(u1p_11) + 2.209012508392e-01*V(u1p_12) + 1.083862483501e-01*V(u1p_13) + 1.289784610271e-01*V(u1p_14)
+ + 1.599046289921e-01*V(u1p_15) + 1.521005928516e-01*V(u1p_16) + -4.721339046955e-02*V(u1p_17) + 5.895599722862e-02*V(u1p_18)
+ + 8.082774281502e-02*V(u1p_19) + 6.992545723915e-02*V(u1m_0) + -4.322490096092e-02*V(u1m_1) + 1.052170991898e-03*V(u1m_2)
+ + -1.664206534624e-01*V(u1m_3) + -4.050457477570e-02*V(u1m_4) + 1.649064421654e-01*V(u1m_5) + -1.753352582455e-02*V(u1m_6)
+ + 1.747005283833e-01*V(u1m_7) + 1.718393862247e-01*V(u1m_8) + 1.166446208954e-01*V(u1m_9) + -3.587155044079e-02*V(u1m_10)
+ + 1.965202689171e-01*V(u1m_11) + 1.127580404282e-01*V(u1m_12) + -2.177745997906e-01*V(u1m_13) + -2.144685536623e-01*V(u1m_14)
+ + -1.371018588543e-01*V(u1m_15) + -1.702023148537e-01*V(u1m_16) + -1.338601708412e-01*V(u1m_17) + 9.209856390953e-02*V(u1m_18)
+ + -1.849099546671e-01*V(u1m_19))
B_u2c_15 u2c_15 0 V = tanh_psi(0.0 + -1.749980449677e-02*(V(u1p_0) + (-1)*V(u1m_0)) + 1.978994607925e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + -8.177617192268e-02*(V(u1p_2) + (-1)*V(u1m_2)) + -1.047352403402e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.471031010151e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + -1.558449864388e-01*(V(u1p_5) + (-1)*V(u1m_5)) + 1.960289180279e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + 5.721926689148e-02*(V(u1p_7) + (-1)*V(u1m_7)) + -5.987411737442e-02*(V(u1p_8) + (-1)*V(u1m_8)) + 8.335164189339e-02*(V(u1p_9)
+ + (-1)*V(u1m_9)) + 4.757893085480e-02*(V(u1p_10) + (-1)*V(u1m_10)) + 7.439351081848e-02*(V(u1p_11) + (-1)*V(u1m_11))
+ + 1.745983064175e-01*(V(u1p_12) + (-1)*V(u1m_12)) + -1.365398466587e-01*(V(u1p_13) + (-1)*V(u1m_13))
+ + -6.879597902298e-03*(V(u1p_14) + (-1)*V(u1m_14)) + 1.736892759800e-01*(V(u1p_15) + (-1)*V(u1m_15)) + 4.402264952660e-03*(V(u1p_16)
+ + (-1)*V(u1m_16)) + 1.494552195072e-01*(V(u1p_17) + (-1)*V(u1m_17)) + 1.992309391499e-01*(V(u1p_18) + (-1)*V(u1m_18))
+ + -8.549882471561e-02*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_16 u2a_16 0 V = tanh_psi(-2.794786989689e-01 + 2.014596164227e-01*V(u1p_0) + -1.943699568510e-01*V(u1p_1) + 6.095120310783e-02*V(u1p_2)
+ + -1.621797084808e-01*V(u1p_3) + -2.113026529551e-01*V(u1p_4) + 7.159736752510e-02*V(u1p_5) + 1.140315830708e-01*V(u1p_6)
+ + 1.356390416622e-01*V(u1p_7) + 2.167009711266e-01*V(u1p_8) + -1.611793041229e-02*V(u1p_9) + 1.084207296371e-01*V(u1p_10)
+ + 1.484425365925e-01*V(u1p_11) + 1.042977869511e-01*V(u1p_12) + -4.885451495647e-02*V(u1p_13) + -1.832370162010e-01*V(u1p_14)
+ + -2.334567904472e-02*V(u1p_15) + 3.668826818466e-02*V(u1p_16) + -1.235848963261e-01*V(u1p_17) + -2.056284099817e-01*V(u1p_18)
+ + 1.578457653522e-01*V(u1p_19) + 7.155209779739e-02*V(u1m_0) + -1.515113115311e-01*V(u1m_1) + 1.372869312763e-01*V(u1m_2)
+ + -1.112090498209e-01*V(u1m_3) + -1.803622543812e-01*V(u1m_4) + 1.184909939766e-01*V(u1m_5) + 1.699641346931e-01*V(u1m_6)
+ + -1.886258274317e-01*V(u1m_7) + 2.107747793198e-01*V(u1m_8) + -1.250622272491e-01*V(u1m_9) + 2.023901343346e-01*V(u1m_10)
+ + -8.906297385693e-02*V(u1m_11) + 6.019017100334e-02*V(u1m_12) + 1.388478875160e-01*V(u1m_13) + 1.091820895672e-01*V(u1m_14)
+ + -2.975162863731e-02*V(u1m_15) + 3.984040021896e-02*V(u1m_16) + 1.357204020023e-01*V(u1m_17) + 9.772652387619e-02*V(u1m_18)
+ + 4.743045568466e-02*V(u1m_19))
B_u2b_16 u2b_16 0 V = tanh_psi(-2.794786989689e-01 + 7.155209779739e-02*V(u1p_0) + -1.515113115311e-01*V(u1p_1) + 1.372869312763e-01*V(u1p_2)
+ + -1.112090498209e-01*V(u1p_3) + -1.803622543812e-01*V(u1p_4) + 1.184909939766e-01*V(u1p_5) + 1.699641346931e-01*V(u1p_6)
+ + -1.886258274317e-01*V(u1p_7) + 2.107747793198e-01*V(u1p_8) + -1.250622272491e-01*V(u1p_9) + 2.023901343346e-01*V(u1p_10)
+ + -8.906297385693e-02*V(u1p_11) + 6.019017100334e-02*V(u1p_12) + 1.388478875160e-01*V(u1p_13) + 1.091820895672e-01*V(u1p_14)
+ + -2.975162863731e-02*V(u1p_15) + 3.984040021896e-02*V(u1p_16) + 1.357204020023e-01*V(u1p_17) + 9.772652387619e-02*V(u1p_18)
+ + 4.743045568466e-02*V(u1p_19) + 2.014596164227e-01*V(u1m_0) + -1.943699568510e-01*V(u1m_1) + 6.095120310783e-02*V(u1m_2)
+ + -1.621797084808e-01*V(u1m_3) + -2.113026529551e-01*V(u1m_4) + 7.159736752510e-02*V(u1m_5) + 1.140315830708e-01*V(u1m_6)
+ + 1.356390416622e-01*V(u1m_7) + 2.167009711266e-01*V(u1m_8) + -1.611793041229e-02*V(u1m_9) + 1.084207296371e-01*V(u1m_10)
+ + 1.484425365925e-01*V(u1m_11) + 1.042977869511e-01*V(u1m_12) + -4.885451495647e-02*V(u1m_13) + -1.832370162010e-01*V(u1m_14)
+ + -2.334567904472e-02*V(u1m_15) + 3.668826818466e-02*V(u1m_16) + -1.235848963261e-01*V(u1m_17) + -2.056284099817e-01*V(u1m_18)
+ + 1.578457653522e-01*V(u1m_19))
B_u2c_16 u2c_16 0 V = tanh_psi(0.0 + 1.339041590691e-01*(V(u1p_0) + (-1)*V(u1m_0)) + -1.041449680924e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + -1.440360248089e-01*(V(u1p_2) + (-1)*V(u1m_2)) + 1.232913434505e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.580290496349e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 7.714912295341e-02*(V(u1p_5) + (-1)*V(u1m_5)) + 8.195084333420e-02*(V(u1p_6) + (-1)*V(u1m_6))
+ + 6.656044721603e-02*(V(u1p_7) + (-1)*V(u1m_7)) + -1.613650768995e-01*(V(u1p_8) + (-1)*V(u1m_8)) + 4.389438033104e-02*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -8.010084927082e-02*(V(u1p_10) + (-1)*V(u1m_10)) + -1.748838722706e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + -7.807104289532e-02*(V(u1p_12) + (-1)*V(u1m_12)) + 1.518179476261e-01*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.614783853292e-01*(V(u1p_14) + (-1)*V(u1m_14)) + 2.194254994392e-01*(V(u1p_15) + (-1)*V(u1m_15)) + 5.701139569283e-02*(V(u1p_16)
+ + (-1)*V(u1m_16)) + -5.547197163105e-02*(V(u1p_17) + (-1)*V(u1m_17)) + -1.687419414520e-01*(V(u1p_18) + (-1)*V(u1m_18))
+ + 1.888367533684e-02*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_17 u2a_17 0 V = tanh_psi(3.193357586861e-02 + -1.958933770657e-01*V(u1p_0) + 5.917075276375e-02*V(u1p_1) + -1.933836489916e-01*V(u1p_2)
+ + -1.340535134077e-01*V(u1p_3) + -2.018417865038e-01*V(u1p_4) + -3.184944391251e-03*V(u1p_5) + -3.276206552982e-02*V(u1p_6)
+ + 4.089367389679e-02*V(u1p_7) + 7.837733626366e-02*V(u1p_8) + 2.862355113029e-02*V(u1p_9) + -1.791701316833e-01*V(u1p_10)
+ + 1.079573631287e-01*V(u1p_11) + -2.020634710789e-02*V(u1p_12) + -1.446799337864e-01*V(u1p_13) + -1.411480903625e-01*V(u1p_14)
+ + -1.080885604024e-01*V(u1p_15) + -1.616009175777e-01*V(u1p_16) + -5.314858257771e-02*V(u1p_17) + -1.978557556868e-01*V(u1p_18)
+ + 1.767451763153e-01*V(u1p_19) + -2.015399634838e-01*V(u1m_0) + 9.539362788200e-02*V(u1m_1) + 2.242186665535e-02*V(u1m_2)
+ + 9.555804729462e-02*V(u1m_3) + -9.415440261364e-02*V(u1m_4) + -2.050692439079e-01*V(u1m_5) + 5.617517232895e-02*V(u1m_6)
+ + 1.918563544750e-01*V(u1m_7) + 1.069269180298e-01*V(u1m_8) + -2.422156929970e-02*V(u1m_9) + 6.522825360298e-02*V(u1m_10)
+ + -2.222283929586e-01*V(u1m_11) + -2.228680551052e-01*V(u1m_12) + 4.611140489578e-02*V(u1m_13) + 1.434774696827e-01*V(u1m_14)
+ + -9.112218022346e-02*V(u1m_15) + 1.509619653225e-01*V(u1m_16) + 2.196224331856e-01*V(u1m_17) + -1.243853792548e-01*V(u1m_18)
+ + 8.152455091476e-02*V(u1m_19))
B_u2b_17 u2b_17 0 V = tanh_psi(3.193357586861e-02 + -2.015399634838e-01*V(u1p_0) + 9.539362788200e-02*V(u1p_1) + 2.242186665535e-02*V(u1p_2)
+ + 9.555804729462e-02*V(u1p_3) + -9.415440261364e-02*V(u1p_4) + -2.050692439079e-01*V(u1p_5) + 5.617517232895e-02*V(u1p_6)
+ + 1.918563544750e-01*V(u1p_7) + 1.069269180298e-01*V(u1p_8) + -2.422156929970e-02*V(u1p_9) + 6.522825360298e-02*V(u1p_10)
+ + -2.222283929586e-01*V(u1p_11) + -2.228680551052e-01*V(u1p_12) + 4.611140489578e-02*V(u1p_13) + 1.434774696827e-01*V(u1p_14)
+ + -9.112218022346e-02*V(u1p_15) + 1.509619653225e-01*V(u1p_16) + 2.196224331856e-01*V(u1p_17) + -1.243853792548e-01*V(u1p_18)
+ + 8.152455091476e-02*V(u1p_19) + -1.958933770657e-01*V(u1m_0) + 5.917075276375e-02*V(u1m_1) + -1.933836489916e-01*V(u1m_2)
+ + -1.340535134077e-01*V(u1m_3) + -2.018417865038e-01*V(u1m_4) + -3.184944391251e-03*V(u1m_5) + -3.276206552982e-02*V(u1m_6)
+ + 4.089367389679e-02*V(u1m_7) + 7.837733626366e-02*V(u1m_8) + 2.862355113029e-02*V(u1m_9) + -1.791701316833e-01*V(u1m_10)
+ + 1.079573631287e-01*V(u1m_11) + -2.020634710789e-02*V(u1m_12) + -1.446799337864e-01*V(u1m_13) + -1.411480903625e-01*V(u1m_14)
+ + -1.080885604024e-01*V(u1m_15) + -1.616009175777e-01*V(u1m_16) + -5.314858257771e-02*V(u1m_17) + -1.978557556868e-01*V(u1m_18)
+ + 1.767451763153e-01*V(u1m_19))
B_u2c_17 u2c_17 0 V = tanh_psi(0.0 + -7.268525660038e-02*(V(u1p_0) + (-1)*V(u1m_0)) + -7.576332986355e-02*(V(u1p_1) + (-1)*V(u1m_1))
+ + -5.553622543812e-02*(V(u1p_2) + (-1)*V(u1m_2)) + -1.837760806084e-01*(V(u1p_3) + (-1)*V(u1m_3)) + -1.671228408813e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + -1.675423830748e-01*(V(u1p_5) + (-1)*V(u1m_5)) + 1.453271508217e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + 3.582930564880e-02*(V(u1p_7) + (-1)*V(u1m_7)) + -2.024227827787e-01*(V(u1p_8) + (-1)*V(u1m_8)) + 1.987786591053e-02*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -8.299641311169e-02*(V(u1p_10) + (-1)*V(u1m_10)) + 1.346732378006e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + 4.822099208832e-02*(V(u1p_12) + (-1)*V(u1m_12)) + -5.598808825016e-02*(V(u1p_13) + (-1)*V(u1m_13)) + 9.076306223869e-02*(V(u1p_14)
+ + (-1)*V(u1m_14)) + -1.140681728721e-01*(V(u1p_15) + (-1)*V(u1m_15)) + 2.075709700584e-01*(V(u1p_16) + (-1)*V(u1m_16))
+ + -7.324564456940e-02*(V(u1p_17) + (-1)*V(u1m_17)) + -9.732022881508e-02*(V(u1p_18) + (-1)*V(u1m_18))
+ + 6.541019678116e-02*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_18 u2a_18 0 V = tanh_psi(-1.348202228546e-01 + -1.510499715805e-01*V(u1p_0) + -8.688603341579e-02*V(u1p_1) + 4.544639587402e-02*V(u1p_2)
+ + 3.923040628433e-02*V(u1p_3) + 2.709829807281e-02*V(u1p_4) + 1.098240315914e-01*V(u1p_5) + -1.841200292110e-01*V(u1p_6)
+ + -1.996058076620e-01*V(u1p_7) + -1.899617612362e-01*V(u1p_8) + -1.599600017071e-01*V(u1p_9) + -1.321371346712e-01*V(u1p_10)
+ + 1.651942729950e-04*V(u1p_11) + -1.145223379135e-01*V(u1p_12) + -2.173388749361e-01*V(u1p_13) + -9.636746346951e-02*V(u1p_14)
+ + 1.384453177452e-01*V(u1p_15) + 1.648893058300e-01*V(u1p_16) + 1.017972528934e-01*V(u1p_17) + 1.190632879734e-01*V(u1p_18)
+ + 1.405905187130e-02*V(u1p_19) + -1.256070733070e-01*V(u1m_0) + -3.158262372017e-02*V(u1m_1) + -5.629602074623e-02*V(u1m_2)
+ + 9.639292955399e-02*V(u1m_3) + -1.689479351044e-01*V(u1m_4) + 1.216866075993e-02*V(u1m_5) + 6.448507308960e-02*V(u1m_6)
+ + -5.781096220016e-02*V(u1m_7) + 7.701396942139e-03*V(u1m_8) + 1.839290261269e-01*V(u1m_9) + 7.066917419434e-02*V(u1m_10)
+ + -1.531242430210e-01*V(u1m_11) + 3.123182058334e-02*V(u1m_12) + 1.887734830379e-01*V(u1m_13) + -1.982637643814e-01*V(u1m_14)
+ + 1.365461945534e-01*V(u1m_15) + 1.527875363827e-01*V(u1m_16) + -5.406825244427e-02*V(u1m_17) + 1.088936924934e-01*V(u1m_18)
+ + -1.864776462317e-01*V(u1m_19))
B_u2b_18 u2b_18 0 V = tanh_psi(-1.348202228546e-01 + -1.256070733070e-01*V(u1p_0) + -3.158262372017e-02*V(u1p_1) + -5.629602074623e-02*V(u1p_2)
+ + 9.639292955399e-02*V(u1p_3) + -1.689479351044e-01*V(u1p_4) + 1.216866075993e-02*V(u1p_5) + 6.448507308960e-02*V(u1p_6)
+ + -5.781096220016e-02*V(u1p_7) + 7.701396942139e-03*V(u1p_8) + 1.839290261269e-01*V(u1p_9) + 7.066917419434e-02*V(u1p_10)
+ + -1.531242430210e-01*V(u1p_11) + 3.123182058334e-02*V(u1p_12) + 1.887734830379e-01*V(u1p_13) + -1.982637643814e-01*V(u1p_14)
+ + 1.365461945534e-01*V(u1p_15) + 1.527875363827e-01*V(u1p_16) + -5.406825244427e-02*V(u1p_17) + 1.088936924934e-01*V(u1p_18)
+ + -1.864776462317e-01*V(u1p_19) + -1.510499715805e-01*V(u1m_0) + -8.688603341579e-02*V(u1m_1) + 4.544639587402e-02*V(u1m_2)
+ + 3.923040628433e-02*V(u1m_3) + 2.709829807281e-02*V(u1m_4) + 1.098240315914e-01*V(u1m_5) + -1.841200292110e-01*V(u1m_6)
+ + -1.996058076620e-01*V(u1m_7) + -1.899617612362e-01*V(u1m_8) + -1.599600017071e-01*V(u1m_9) + -1.321371346712e-01*V(u1m_10)
+ + 1.651942729950e-04*V(u1m_11) + -1.145223379135e-01*V(u1m_12) + -2.173388749361e-01*V(u1m_13) + -9.636746346951e-02*V(u1m_14)
+ + 1.384453177452e-01*V(u1m_15) + 1.648893058300e-01*V(u1m_16) + 1.017972528934e-01*V(u1m_17) + 1.190632879734e-01*V(u1m_18)
+ + 1.405905187130e-02*V(u1m_19))
B_u2c_18 u2c_18 0 V = tanh_psi(0.0 + -9.784409403801e-02*(V(u1p_0) + (-1)*V(u1m_0)) + -1.843700557947e-01*(V(u1p_1) + (-1)*V(u1m_1))
+ + 7.982409000397e-02*(V(u1p_2) + (-1)*V(u1m_2)) + 3.801620006561e-02*(V(u1p_3) + (-1)*V(u1m_3)) + -8.871486783028e-02*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 6.562617421150e-02*(V(u1p_5) + (-1)*V(u1m_5)) + -1.628329157829e-01*(V(u1p_6) + (-1)*V(u1m_6))
+ + 9.373578429222e-02*(V(u1p_7) + (-1)*V(u1m_7)) + 2.647405862808e-02*(V(u1p_8) + (-1)*V(u1m_8)) + 1.577903926373e-01*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -7.590055465698e-02*(V(u1p_10) + (-1)*V(u1m_10)) + 1.267231702805e-01*(V(u1p_11) + (-1)*V(u1m_11))
+ + 1.215599477291e-01*(V(u1p_12) + (-1)*V(u1m_12)) + -2.044198065996e-01*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.881833374500e-01*(V(u1p_14) + (-1)*V(u1m_14)) + 1.733478009701e-01*(V(u1p_15) + (-1)*V(u1m_15)) + 2.066827416420e-01*(V(u1p_16)
+ + (-1)*V(u1m_16)) + 1.654627025127e-01*(V(u1p_17) + (-1)*V(u1m_17)) + -2.007442861795e-01*(V(u1p_18) + (-1)*V(u1m_18))
+ + -1.097744479775e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u2a_19 u2a_19 0 V = tanh_psi(1.554517447948e-02 + 2.355201542377e-02*V(u1p_0) + -1.610064655542e-01*V(u1p_1) + -1.074399426579e-01*V(u1p_2)
+ + -1.937505006790e-01*V(u1p_3) + 3.720268607140e-03*V(u1p_4) + -3.375647962093e-02*V(u1p_5) + -2.033351957798e-01*V(u1p_6)
+ + -1.069766357541e-01*V(u1p_7) + 3.824263811111e-03*V(u1p_8) + -1.015354245901e-01*V(u1p_9) + 2.095807194710e-01*V(u1p_10)
+ + -1.610046625137e-01*V(u1p_11) + -1.260014772415e-01*V(u1p_12) + 4.950308799744e-02*V(u1p_13) + 2.194127440453e-02*V(u1p_14)
+ + 1.529865562916e-01*V(u1p_15) + 3.488963842392e-02*V(u1p_16) + 3.055429458618e-02*V(u1p_17) + -2.082148194313e-01*V(u1p_18)
+ + -1.498776674271e-02*V(u1p_19) + -4.952606558800e-02*V(u1m_0) + 1.199741363525e-01*V(u1m_1) + -1.658463180065e-01*V(u1m_2)
+ + -1.895303428173e-01*V(u1m_3) + 7.235679030418e-02*V(u1m_4) + -1.834631711245e-01*V(u1m_5) + -1.455379128456e-01*V(u1m_6)
+ + 1.308380067348e-02*V(u1m_7) + -4.111433029175e-02*V(u1m_8) + -4.774302244186e-03*V(u1m_9) + 2.104663848877e-01*V(u1m_10)
+ + 1.887737512589e-01*V(u1m_11) + 1.236221790314e-01*V(u1m_12) + -7.567451894283e-02*V(u1m_13) + -2.881194651127e-02*V(u1m_14)
+ + -3.341042995453e-02*V(u1m_15) + 1.930991113186e-01*V(u1m_16) + 2.084315121174e-01*V(u1m_17) + -6.355136632919e-03*V(u1m_18)
+ + -1.057006642222e-01*V(u1m_19))
B_u2b_19 u2b_19 0 V = tanh_psi(1.554517447948e-02 + -4.952606558800e-02*V(u1p_0) + 1.199741363525e-01*V(u1p_1) + -1.658463180065e-01*V(u1p_2)
+ + -1.895303428173e-01*V(u1p_3) + 7.235679030418e-02*V(u1p_4) + -1.834631711245e-01*V(u1p_5) + -1.455379128456e-01*V(u1p_6)
+ + 1.308380067348e-02*V(u1p_7) + -4.111433029175e-02*V(u1p_8) + -4.774302244186e-03*V(u1p_9) + 2.104663848877e-01*V(u1p_10)
+ + 1.887737512589e-01*V(u1p_11) + 1.236221790314e-01*V(u1p_12) + -7.567451894283e-02*V(u1p_13) + -2.881194651127e-02*V(u1p_14)
+ + -3.341042995453e-02*V(u1p_15) + 1.930991113186e-01*V(u1p_16) + 2.084315121174e-01*V(u1p_17) + -6.355136632919e-03*V(u1p_18)
+ + -1.057006642222e-01*V(u1p_19) + 2.355201542377e-02*V(u1m_0) + -1.610064655542e-01*V(u1m_1) + -1.074399426579e-01*V(u1m_2)
+ + -1.937505006790e-01*V(u1m_3) + 3.720268607140e-03*V(u1m_4) + -3.375647962093e-02*V(u1m_5) + -2.033351957798e-01*V(u1m_6)
+ + -1.069766357541e-01*V(u1m_7) + 3.824263811111e-03*V(u1m_8) + -1.015354245901e-01*V(u1m_9) + 2.095807194710e-01*V(u1m_10)
+ + -1.610046625137e-01*V(u1m_11) + -1.260014772415e-01*V(u1m_12) + 4.950308799744e-02*V(u1m_13) + 2.194127440453e-02*V(u1m_14)
+ + 1.529865562916e-01*V(u1m_15) + 3.488963842392e-02*V(u1m_16) + 3.055429458618e-02*V(u1m_17) + -2.082148194313e-01*V(u1m_18)
+ + -1.498776674271e-02*V(u1m_19))
B_u2c_19 u2c_19 0 V = tanh_psi(0.0 + -8.809636533260e-02*(V(u1p_0) + (-1)*V(u1m_0)) + 3.209826350212e-02*(V(u1p_1) + (-1)*V(u1m_1))
+ + -1.081880182028e-01*(V(u1p_2) + (-1)*V(u1m_2)) + -1.023733019829e-01*(V(u1p_3) + (-1)*V(u1m_3)) + 1.175428926945e-01*(V(u1p_4)
+ + (-1)*V(u1m_4)) + 6.564071774483e-02*(V(u1p_5) + (-1)*V(u1m_5)) + 4.910796880722e-02*(V(u1p_6) + (-1)*V(u1m_6))
+ + -6.658463180065e-02*(V(u1p_7) + (-1)*V(u1m_7)) + 2.925604581833e-02*(V(u1p_8) + (-1)*V(u1m_8)) + -1.088033616543e-02*(V(u1p_9)
+ + (-1)*V(u1m_9)) + -6.669023633003e-02*(V(u1p_10) + (-1)*V(u1m_10)) + 7.468175888062e-02*(V(u1p_11) + (-1)*V(u1m_11))
+ + -2.015954405069e-01*(V(u1p_12) + (-1)*V(u1m_12)) + -9.069392085075e-02*(V(u1p_13) + (-1)*V(u1m_13))
+ + -1.099647730589e-01*(V(u1p_14) + (-1)*V(u1m_14)) + -8.496570587158e-02*(V(u1p_15) + (-1)*V(u1m_15))
+ + 1.965708434582e-01*(V(u1p_16) + (-1)*V(u1m_16)) + 2.203918099403e-01*(V(u1p_17) + (-1)*V(u1m_17)) + -1.745047718287e-01*(V(u1p_18)
+ + (-1)*V(u1m_18)) + 1.807030737400e-01*(V(u1p_19) + (-1)*V(u1m_19)))
B_u3_0 u3_0 0 V = tanh_psi(0.0 + 3.581413626671e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -1.671868860722e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 2.136018276215e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 1.235789060593e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -1.858746111393e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -2.313661575317e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 8.581098914146e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 5.254730582237e-03*(V(u2a_7) + (-1)*V(u2b_7)) + -5.668528378010e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -1.063790321350e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 7.425913214684e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 4.687356948853e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 1.375851631165e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 1.938866376877e-01*(V(u2a_13) + (-1)*V(u2b_13)) + -1.639090925455e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + 4.938572645187e-02*(V(u2a_15) + (-1)*V(u2b_15)) + -1.795876026154e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + 2.030852437019e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -9.403607249260e-02*(V(u2a_18) + (-1)*V(u2b_18))
+ + -1.380571722984e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 1.836506128311e-01*V(u2c_0) + -2.347354590893e-02*V(u2c_1)
+ + -1.267249882221e-01*V(u2c_2) + -9.103685617447e-03*V(u2c_3) + 5.128982663155e-02*V(u2c_4) + -6.207972764969e-03*V(u2c_5)
+ + -2.108627408743e-01*V(u2c_6) + -1.894810199738e-01*V(u2c_7) + 9.630128741264e-02*V(u2c_8) + -1.100086197257e-01*V(u2c_9)
+ + -2.855753898621e-02*V(u2c_10) + 1.757260560989e-01*V(u2c_11) + -1.867900788784e-01*V(u2c_12) + 1.483039557934e-02*V(u2c_13)
+ + -2.141357511282e-01*V(u2c_14) + 7.116135954857e-02*V(u2c_15) + -1.259966492653e-01*V(u2c_16) + -6.203903257847e-02*V(u2c_17)
+ + -8.521883189678e-02*V(u2c_18) + 4.999512434006e-02*V(u2c_19))
B_u3_1 u3_1 0 V = tanh_psi(0.0 + 1.282262802124e-02*(V(u2a_0) + (-1)*V(u2b_0)) + 6.307181715965e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + 8.671581745148e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 8.771350979805e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -1.295440644026e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 1.873581409454e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 1.099877655506e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -3.994661569595e-02*(V(u2a_7) + (-1)*V(u2b_7)) + -1.774360239506e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -8.044023811817e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.040001735091e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -1.864158213139e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.907164007425e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 1.524982750416e-01*(V(u2a_13) + (-1)*V(u2b_13)) + 1.488081514835e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.360446810722e-01*(V(u2a_15) + (-1)*V(u2b_15)) + -7.682372629642e-02*(V(u2a_16) + (-1)*V(u2b_16))
+ + 1.681885123253e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 1.852299273014e-01*(V(u2a_18) + (-1)*V(u2b_18)) + 1.017300784588e-01*(V(u2a_19)
+ + (-1)*V(u2b_19)) + -2.136035114527e-01*V(u2c_0) + 1.467714011669e-01*V(u2c_1) + 1.641088426113e-01*V(u2c_2)
+ + -2.168142795563e-01*V(u2c_3) + -4.645872116089e-02*V(u2c_4) + -2.087536901236e-01*V(u2c_5) + 2.898311614990e-02*V(u2c_6)
+ + -1.326712667942e-01*V(u2c_7) + 1.002067029476e-01*V(u2c_8) + 1.586858928204e-02*V(u2c_9) + -1.387287676334e-02*V(u2c_10)
+ + 9.530404210091e-02*V(u2c_11) + 4.270529747009e-02*V(u2c_12) + -1.378460526466e-01*V(u2c_13) + 2.062414586544e-01*V(u2c_14)
+ + 1.245246231556e-01*V(u2c_15) + -2.201129645109e-01*V(u2c_16) + -1.105565354228e-01*V(u2c_17) + -7.147920131683e-02*V(u2c_18)
+ + -3.514513373375e-03*V(u2c_19))
B_u3_2 u3_2 0 V = tanh_psi(0.0 + 1.366804838181e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 2.115304172039e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 7.103836536407e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -2.329559624195e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -1.208642572165e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.711836010218e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 1.390978991985e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -5.304031074047e-02*(V(u2a_7) + (-1)*V(u2b_7)) + -2.072483301163e-03*(V(u2a_8) + (-1)*V(u2b_8)) + -1.019688248634e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 2.889606356621e-02*(V(u2a_10) + (-1)*V(u2b_10)) + -4.045635461807e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + -7.096193730831e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 9.499433636665e-02*(V(u2a_13) + (-1)*V(u2b_13)) + 1.545773446560e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -2.045038938522e-01*(V(u2a_15) + (-1)*V(u2b_15)) + -1.504815071821e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + 2.464517951012e-02*(V(u2a_17) + (-1)*V(u2b_17)) + -8.850732445717e-02*(V(u2a_18) + (-1)*V(u2b_18)) + 2.104779779911e-01*(V(u2a_19)
+ + (-1)*V(u2b_19)) + 1.299339532852e-02*V(u2c_0) + -1.498106718063e-01*V(u2c_1) + 5.505970120430e-02*V(u2c_2)
+ + 5.191698670387e-02*V(u2c_3) + 6.341460347176e-02*V(u2c_4) + -1.676522642374e-01*V(u2c_5) + -6.621426343918e-02*V(u2c_6)
+ + -1.651305556297e-01*V(u2c_7) + 1.011165976524e-02*V(u2c_8) + -1.716871857643e-01*V(u2c_9) + 1.680388748646e-01*V(u2c_10)
+ + 9.681606292725e-02*V(u2c_11) + 1.087377965450e-02*V(u2c_12) + 1.446350812912e-01*V(u2c_13) + 6.470182538033e-02*V(u2c_14)
+ + 4.891765117645e-02*V(u2c_15) + 1.770831346512e-01*V(u2c_16) + 2.005577683449e-01*V(u2c_17) + -1.326081752777e-01*V(u2c_18)
+ + 1.450249552727e-01*V(u2c_19))
B_u3_3 u3_3 0 V = tanh_psi(0.0 + 2.065036594868e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 1.848659217358e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 7.661539316177e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 1.782298982143e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 5.861249566078e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.513718068600e-01*(V(u2a_5) + (-1)*V(u2b_5)) + -6.231756508350e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.427075266838e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 1.393203437328e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 2.118546366692e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -2.175751775503e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 9.209603071213e-03*(V(u2a_11) + (-1)*V(u2b_11))
+ + -8.032332360744e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 1.215083301067e-01*(V(u2a_13) + (-1)*V(u2b_13))
+ + -2.145927697420e-01*(V(u2a_14) + (-1)*V(u2b_14)) + 1.473736763000e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 1.710014045238e-01*(V(u2a_16)
+ + (-1)*V(u2b_16)) + -1.195135116577e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -2.096483558416e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + 8.702334761620e-02*(V(u2a_19) + (-1)*V(u2b_19)) + 1.412655413151e-01*V(u2c_0) + -1.471903026104e-01*V(u2c_1)
+ + 1.431657671928e-01*V(u2c_2) + -1.153471767902e-01*V(u2c_3) + -2.806845307350e-02*V(u2c_4) + 3.897437453270e-02*V(u2c_5)
+ + -7.880933582783e-02*V(u2c_6) + 2.150090038776e-02*V(u2c_7) + -1.567250490189e-02*V(u2c_8) + -1.132466867566e-01*V(u2c_9)
+ + 1.138149797916e-01*V(u2c_10) + 2.016029357910e-01*V(u2c_11) + 9.389585256577e-02*V(u2c_12) + 1.464727520943e-01*V(u2c_13)
+ + -1.855262815952e-01*V(u2c_14) + -1.096018254757e-01*V(u2c_15) + 7.098054885864e-02*V(u2c_16) + 1.841973960400e-01*V(u2c_17)
+ + -1.791357994080e-03*V(u2c_18) + -1.760219633579e-01*V(u2c_19))
B_u3_4 u3_4 0 V = tanh_psi(0.0 + -1.633770167828e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 1.736180186272e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 8.505770564079e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -1.750776916742e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -8.036527037621e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -2.683937549591e-03*(V(u2a_5) + (-1)*V(u2b_5)) + -4.934200644493e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.755826175213e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 3.980606794357e-02*(V(u2a_8) + (-1)*V(u2b_8)) + 1.534378826618e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 9.241196513176e-02*(V(u2a_10) + (-1)*V(u2b_10)) + -9.471563994884e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + -9.754467010498e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 1.932130157948e-01*(V(u2a_13) + (-1)*V(u2b_13))
+ + -4.086965322495e-02*(V(u2a_14) + (-1)*V(u2b_14)) + 3.085634112358e-02*(V(u2a_15) + (-1)*V(u2b_15))
+ + -2.192614078522e-01*(V(u2a_16) + (-1)*V(u2b_16)) + -7.184934616089e-02*(V(u2a_17) + (-1)*V(u2b_17))
+ + -1.908372342587e-01*(V(u2a_18) + (-1)*V(u2b_18)) + -2.693419158459e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -8.384883403778e-04*V(u2c_0)
+ + -9.039899706841e-02*V(u2c_1) + -6.343244016171e-02*V(u2c_2) + -1.346930861473e-02*V(u2c_3) + -1.087439805269e-01*V(u2c_4)
+ + -9.306097030640e-02*V(u2c_5) + -1.637234836817e-01*V(u2c_6) + -1.162412464619e-01*V(u2c_7) + 2.090243995190e-02*V(u2c_8)
+ + 3.229424357414e-03*V(u2c_9) + -6.608031690121e-02*V(u2c_10) + 1.796954870224e-01*V(u2c_11) + 3.597718477249e-02*V(u2c_12)
+ + -1.955221891403e-01*V(u2c_13) + 3.367203474045e-02*V(u2c_14) + -3.617966175079e-02*V(u2c_15) + -9.748555719852e-02*V(u2c_16)
+ + 2.113394737244e-01*V(u2c_17) + -3.205849230289e-02*V(u2c_18) + -1.987459957600e-01*V(u2c_19))
B_u3_5 u3_5 0 V = tanh_psi(0.0 + 1.438190042973e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -2.195118516684e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 3.624573349953e-03*(V(u2a_2) + (-1)*V(u2b_2)) + 2.158662676811e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -5.397678911686e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 1.521714627743e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 5.490052700043e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 6.400993466377e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 2.051476836205e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.249576807022e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.466932296753e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 4.303067922592e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 1.876716315746e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 1.321406066418e-01*(V(u2a_13) + (-1)*V(u2b_13)) + -2.027423083782e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + 1.218115389347e-01*(V(u2a_15) + (-1)*V(u2b_15)) + -6.004151701927e-02*(V(u2a_16) + (-1)*V(u2b_16))
+ + 1.434950828552e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -2.228233963251e-01*(V(u2a_18) + (-1)*V(u2b_18)) + 1.993253231049e-01*(V(u2a_19)
+ + (-1)*V(u2b_19)) + 7.780426740646e-02*V(u2c_0) + 2.885848283768e-02*V(u2c_1) + 3.412380814552e-02*V(u2c_2)
+ + -7.086968421936e-02*V(u2c_3) + 1.343605518341e-01*V(u2c_4) + -4.395431280136e-02*V(u2c_5) + -4.382118582726e-03*V(u2c_6)
+ + 1.945739686489e-01*V(u2c_7) + -5.285139381886e-02*V(u2c_8) + 1.830069422722e-01*V(u2c_9) + 1.111581921577e-01*V(u2c_10)
+ + 1.647091507912e-01*V(u2c_11) + 5.277267098427e-02*V(u2c_12) + 6.289017200470e-02*V(u2c_13) + 2.180569469929e-01*V(u2c_14)
+ + -1.549292802811e-01*V(u2c_15) + -4.589170217514e-02*V(u2c_16) + -1.070851534605e-01*V(u2c_17) + -1.163186058402e-01*V(u2c_18)
+ + 5.304417014122e-02*V(u2c_19))
B_u3_6 u3_6 0 V = tanh_psi(0.0 + 2.118257582188e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 1.097541749477e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 4.558730125427e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -1.220982670784e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -1.589593142271e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 2.106679677963e-01*(V(u2a_5) + (-1)*V(u2b_5)) + -1.307296156883e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.801293790340e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -1.131062880158e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 2.831286191940e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -3.471601009369e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.991426348686e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.987203210592e-01*(V(u2a_12) + (-1)*V(u2b_12)) + -2.293059229851e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + -5.473797023296e-02*(V(u2a_14) + (-1)*V(u2b_14)) + 1.870133876801e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 7.427930831909e-04*(V(u2a_16)
+ + (-1)*V(u2b_16)) + -1.425924003124e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 5.046710371971e-02*(V(u2a_18) + (-1)*V(u2b_18))
+ + -1.833514273167e-01*(V(u2a_19) + (-1)*V(u2b_19)) + -5.895379185677e-02*V(u2c_0) + 4.808047413826e-02*V(u2c_1)
+ + 2.179310321808e-01*V(u2c_2) + -1.241407543421e-01*V(u2c_3) + -2.009174227715e-01*V(u2c_4) + 9.750211238861e-02*V(u2c_5)
+ + 1.856331527233e-01*V(u2c_6) + -1.384185254574e-01*V(u2c_7) + -1.387429535389e-01*V(u2c_8) + 1.625982522964e-01*V(u2c_9)
+ + -2.008050680161e-03*V(u2c_10) + 1.729249954224e-03*V(u2c_11) + 2.295777201653e-03*V(u2c_12) + 9.028100967407e-02*V(u2c_13)
+ + 1.801240146160e-01*V(u2c_14) + 2.628095448017e-02*V(u2c_15) + 1.885806620121e-01*V(u2c_16) + 7.478690147400e-02*V(u2c_17)
+ + -2.034827321768e-01*V(u2c_18) + -1.799806654453e-01*V(u2c_19))
B_u3_7 u3_7 0 V = tanh_psi(0.0 + -1.105481162667e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 1.051932275295e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -6.081381440163e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 3.785407543182e-02*(V(u2a_3) + (-1)*V(u2b_3)) + 6.817331910133e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 2.186138629913e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 2.533821761608e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + -4.932716488838e-03*(V(u2a_7) + (-1)*V(u2b_7)) + 9.453102946281e-03*(V(u2a_8) + (-1)*V(u2b_8)) + 2.076600790024e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 2.058089375496e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -3.989487886429e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + -9.821021556854e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -6.558838486671e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + 5.449089407921e-02*(V(u2a_14) + (-1)*V(u2b_14)) + 1.992697417736e-01*(V(u2a_15) + (-1)*V(u2b_15)) + -7.349868118763e-02*(V(u2a_16)
+ + (-1)*V(u2b_16)) + -4.503178596497e-02*(V(u2a_17) + (-1)*V(u2b_17)) + 1.612319648266e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + 1.579238772392e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 1.984001994133e-01*V(u2c_0) + 7.188808917999e-02*V(u2c_1)
+ + -1.215032786131e-01*V(u2c_2) + 4.643794894218e-02*V(u2c_3) + -8.022874593735e-02*V(u2c_4) + -2.149877548218e-01*V(u2c_5)
+ + 3.691315650940e-02*V(u2c_6) + 1.374844312668e-01*V(u2c_7) + -7.688991725445e-02*V(u2c_8) + 4.819431900978e-02*V(u2c_9)
+ + 1.130447387695e-01*V(u2c_10) + -1.540574431419e-01*V(u2c_11) + -2.112989127636e-01*V(u2c_12) + 4.900747537613e-02*V(u2c_13)
+ + -1.066899299622e-02*V(u2c_14) + 1.642503738403e-01*V(u2c_15) + 1.618042588234e-03*V(u2c_16) + -1.563730239868e-01*V(u2c_17)
+ + 2.124971449375e-01*V(u2c_18) + 1.428088545799e-01*V(u2c_19))
B_u3_8 u3_8 0 V = tanh_psi(0.0 + 1.377715766430e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 1.391646265984e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.954134702682e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -1.711398065090e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -1.242928281426e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.332964301109e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 1.066260933876e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 2.766135334969e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 2.068463265896e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.787413656712e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.908757239580e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 1.573147177696e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 1.524379253387e-01*(V(u2a_12) + (-1)*V(u2b_12)) + -5.444370210171e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + -1.899962425232e-01*(V(u2a_14) + (-1)*V(u2b_14)) + 2.001167535782e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 4.200902581215e-02*(V(u2a_16)
+ + (-1)*V(u2b_16)) + -1.031430065632e-02*(V(u2a_17) + (-1)*V(u2b_17)) + 3.952404856682e-02*(V(u2a_18) + (-1)*V(u2b_18))
+ + 6.770578026772e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -2.028370201588e-01*V(u2c_0) + -7.110060751438e-02*V(u2c_1)
+ + -1.545901298523e-01*V(u2c_2) + 1.253052055836e-01*V(u2c_3) + 1.681021451950e-01*V(u2c_4) + -1.031967848539e-01*V(u2c_5)
+ + -1.180524751544e-01*V(u2c_6) + -1.659048050642e-01*V(u2c_7) + -2.023943364620e-01*V(u2c_8) + 7.890677452087e-02*V(u2c_9)
+ + -1.470737457275e-01*V(u2c_10) + 6.033474206924e-02*V(u2c_11) + -9.998532384634e-02*V(u2c_12) + -5.311244726181e-02*V(u2c_13)
+ + -3.109769523144e-02*V(u2c_14) + -7.567726075649e-02*V(u2c_15) + -2.007536888123e-01*V(u2c_16) + 1.689581871033e-01*V(u2c_17)
+ + -1.877970397472e-01*V(u2c_18) + 5.150145292282e-02*V(u2c_19))
B_u3_9 u3_9 0 V = tanh_psi(0.0 + -9.340251982212e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -1.134753152728e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -4.584294557571e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -1.888788193464e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -1.077416911721e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -4.544971883297e-02*(V(u2a_5) + (-1)*V(u2b_5)) + -2.169585227966e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.239335313439e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 1.209841072559e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.025087237358e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 2.353642880917e-02*(V(u2a_10) + (-1)*V(u2b_10)) + -7.589308917522e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.033707708120e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 1.885386705399e-01*(V(u2a_13) + (-1)*V(u2b_13)) + 1.489835381508e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.143466234207e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 1.761566102505e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + -6.533819437027e-02*(V(u2a_17) + (-1)*V(u2b_17)) + -2.098176479340e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + -2.367207407951e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -7.612942159176e-02*V(u2c_0) + 2.716061472893e-02*V(u2c_1)
+ + 1.865702271461e-01*V(u2c_2) + -2.346664667130e-03*V(u2c_3) + -3.331755101681e-02*V(u2c_4) + 7.957237958908e-02*V(u2c_5)
+ + -1.193692237139e-01*V(u2c_6) + 8.553627133369e-02*V(u2c_7) + -8.602392673492e-02*V(u2c_8) + -4.309943318367e-02*V(u2c_9)
+ + -1.674249768257e-01*V(u2c_10) + -7.059547305107e-02*V(u2c_11) + 2.014230191708e-01*V(u2c_12) + 1.130757331848e-01*V(u2c_13)
+ + 2.037656903267e-01*V(u2c_14) + 1.538397967815e-01*V(u2c_15) + 3.535553812981e-02*V(u2c_16) + 2.081456482410e-01*V(u2c_17)
+ + -1.932666003704e-01*V(u2c_18) + -9.898222982883e-02*V(u2c_19))
B_u3_10 u3_10 0 V = tanh_psi(0.0 + 3.529185056686e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -7.434234023094e-03*(V(u2a_1) + (-1)*V(u2b_1))
+ + -4.429742693901e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -7.516247034073e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -7.188856601715e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -3.149598836899e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 1.998779475689e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.679920703173e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -1.804606914520e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.764782071114e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -2.109850645065e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -1.677364408970e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.052575856447e-01*(V(u2a_12) + (-1)*V(u2b_12)) + -1.046857088804e-01*(V(u2a_13) + (-1)*V(u2b_13))
+ + 1.561420857906e-01*(V(u2a_14) + (-1)*V(u2b_14)) + 2.504502236843e-02*(V(u2a_15) + (-1)*V(u2b_15)) + -1.156458333135e-01*(V(u2a_16)
+ + (-1)*V(u2b_16)) + -2.052537351847e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -1.454748958349e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + 4.589775204659e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -1.390076875687e-01*V(u2c_0) + -1.280285418034e-01*V(u2c_1)
+ + -1.581203341484e-01*V(u2c_2) + 2.775543928146e-02*V(u2c_3) + -1.171926036477e-01*V(u2c_4) + 7.011795043945e-02*V(u2c_5)
+ + -2.055365294218e-01*V(u2c_6) + 8.357715606689e-02*V(u2c_7) + 5.314990878105e-03*V(u2c_8) + 1.098197698593e-02*V(u2c_9)
+ + -1.279413700104e-01*V(u2c_10) + -1.188112050295e-01*V(u2c_11) + -8.696936070919e-02*V(u2c_12) + 5.319178104401e-03*V(u2c_13)
+ + 2.665483951569e-02*V(u2c_14) + -1.473043262959e-01*V(u2c_15) + 1.467221975327e-01*V(u2c_16) + -2.200708985329e-01*V(u2c_17)
+ + 1.946536600590e-01*V(u2c_18) + -1.279786229134e-03*V(u2c_19))
B_u3_11 u3_11 0 V = tanh_psi(0.0 + 2.143856883049e-02*(V(u2a_0) + (-1)*V(u2b_0)) + 1.053603291512e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 2.024473547935e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -1.473731100559e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -1.729341000319e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.461585462093e-01*(V(u2a_5) + (-1)*V(u2b_5)) + -1.173610985279e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -6.439030170441e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 2.138821780682e-01*(V(u2a_8) + (-1)*V(u2b_8)) + -2.064336687326e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -2.041615247726e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 5.935975909233e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 4.798644781113e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 8.514589071274e-02*(V(u2a_13) + (-1)*V(u2b_13)) + -9.436847269535e-02*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.782064735889e-01*(V(u2a_15) + (-1)*V(u2b_15)) + -1.167095974088e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + -1.478819549084e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 8.907595276833e-02*(V(u2a_18) + (-1)*V(u2b_18))
+ + -7.477049529552e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -1.075368076563e-01*V(u2c_0) + 2.065351307392e-01*V(u2c_1)
+ + 4.608938097954e-02*V(u2c_2) + 2.212541997433e-01*V(u2c_3) + -1.078415662050e-01*V(u2c_4) + 1.838076710701e-01*V(u2c_5)
+ + 1.467843353748e-01*V(u2c_6) + 2.029207348824e-01*V(u2c_7) + -1.768509596586e-01*V(u2c_8) + 2.089583277702e-01*V(u2c_9)
+ + 1.434831917286e-01*V(u2c_10) + -8.198617398739e-02*V(u2c_11) + -5.635444819927e-02*V(u2c_12) + 2.009078860283e-02*V(u2c_13)
+ + 9.625747799873e-02*V(u2c_14) + 1.029258370399e-01*V(u2c_15) + -1.711009740829e-01*V(u2c_16) + -6.919243931770e-02*V(u2c_17)
+ + -2.027457207441e-01*V(u2c_18) + -1.599815487862e-01*V(u2c_19))
B_u3_12 u3_12 0 V = tanh_psi(0.0 + -1.561892777681e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.876276731491e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.340434253216e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 1.995694935322e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 1.627866625786e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 1.629185676575e-02*(V(u2a_5) + (-1)*V(u2b_5)) + -4.802380502224e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 7.918885350227e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 8.739674091339e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -2.111410796642e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 9.873390197754e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.383772492409e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 2.051213085651e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 3.314188122749e-02*(V(u2a_13) + (-1)*V(u2b_13)) + -1.101939901710e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.938863843679e-01*(V(u2a_15) + (-1)*V(u2b_15)) + -1.516590565443e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + 3.956294059753e-02*(V(u2a_17) + (-1)*V(u2b_17)) + 1.007646918297e-01*(V(u2a_18) + (-1)*V(u2b_18)) + -2.271395921707e-02*(V(u2a_19)
+ + (-1)*V(u2b_19)) + 1.737743020058e-01*V(u2c_0) + 8.488613367081e-02*V(u2c_1) + 1.381212472916e-02*V(u2c_2)
+ + 4.100680351257e-03*V(u2c_3) + -1.796469688416e-01*V(u2c_4) + -3.899453580379e-02*V(u2c_5) + -8.158484101295e-02*V(u2c_6)
+ + 1.023476719856e-01*V(u2c_7) + 1.700620353222e-01*V(u2c_8) + 6.264585256577e-02*V(u2c_9) + -7.902738451958e-02*V(u2c_10)
+ + 4.979571700096e-02*V(u2c_11) + -1.818347275257e-01*V(u2c_12) + 1.334338486195e-01*V(u2c_13) + -1.202572733164e-01*V(u2c_14)
+ + -5.916644632816e-02*V(u2c_15) + -1.247307062149e-01*V(u2c_16) + -2.234423011541e-01*V(u2c_17) + -6.753949820995e-02*V(u2c_18)
+ + -1.632064133883e-01*V(u2c_19))
B_u3_13 u3_13 0 V = tanh_psi(0.0 + -1.039023175836e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 1.467765569687e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 2.189241349697e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -1.832161247730e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 2.009128034115e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 1.982500553131e-01*(V(u2a_5) + (-1)*V(u2b_5)) + -1.757530868053e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.585722863674e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 8.953762054443e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -2.109613418579e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -7.004514336586e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.791690587997e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.878447830677e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 1.403995156288e-01*(V(u2a_13) + (-1)*V(u2b_13)) + 8.516651391983e-02*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.261567771435e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 8.522647619247e-02*(V(u2a_16) + (-1)*V(u2b_16))
+ + 8.439925312996e-02*(V(u2a_17) + (-1)*V(u2b_17)) + 7.134974002838e-02*(V(u2a_18) + (-1)*V(u2b_18)) + 8.116418123245e-02*(V(u2a_19)
+ + (-1)*V(u2b_19)) + 6.616786122322e-02*V(u2c_0) + 1.075534820557e-01*V(u2c_1) + -1.585410535336e-01*V(u2c_2)
+ + -1.765756905079e-01*V(u2c_3) + -6.932462751865e-02*V(u2c_4) + -1.356005221605e-01*V(u2c_5) + -1.940474957228e-01*V(u2c_6)
+ + -1.199144721031e-01*V(u2c_7) + 1.515430510044e-01*V(u2c_8) + 1.183111965656e-01*V(u2c_9) + 1.615260839462e-01*V(u2c_10)
+ + 2.269361913204e-02*V(u2c_11) + -1.501348614693e-02*V(u2c_12) + 1.927830874920e-01*V(u2c_13) + 2.866241335869e-02*V(u2c_14)
+ + -2.119240760803e-01*V(u2c_15) + -7.684826850891e-03*V(u2c_16) + -8.902847766876e-02*V(u2c_17) + 6.007778644562e-02*V(u2c_18)
+ + 2.006298899651e-01*V(u2c_19))
B_u3_14 u3_14 0 V = tanh_psi(0.0 + -4.324300587177e-02*(V(u2a_0) + (-1)*V(u2b_0)) + 1.062400341034e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.957662105560e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 1.065388321877e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 1.409965455532e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.885889321566e-01*(V(u2a_5) + (-1)*V(u2b_5)) + -1.883883774281e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.661674678326e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -1.890885233879e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.934647560120e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 1.230212450027e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -6.569495797157e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + -6.753513216972e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -2.285413444042e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + -2.207589149475e-01*(V(u2a_14) + (-1)*V(u2b_14)) + -9.376087784767e-02*(V(u2a_15) + (-1)*V(u2b_15))
+ + 1.111433207989e-01*(V(u2a_16) + (-1)*V(u2b_16)) + 2.071703672409e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 1.141229271889e-01*(V(u2a_18)
+ + (-1)*V(u2b_18)) + -5.449794232845e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -8.184894919395e-02*V(u2c_0) + -2.120547741652e-01*V(u2c_1)
+ + -1.873409450054e-01*V(u2c_2) + -1.960960328579e-01*V(u2c_3) + -2.115752100945e-01*V(u2c_4) + 1.942559480667e-01*V(u2c_5)
+ + -1.013686358929e-01*V(u2c_6) + -2.069874107838e-01*V(u2c_7) + -5.804717540741e-03*V(u2c_8) + 1.075895428658e-01*V(u2c_9)
+ + -5.773162841797e-02*V(u2c_10) + -9.782858192921e-02*V(u2c_11) + 5.829799175262e-02*V(u2c_12) + -3.540730476379e-02*V(u2c_13)
+ + 7.827800512314e-02*V(u2c_14) + 1.934243738651e-01*V(u2c_15) + -7.038494944572e-02*V(u2c_16) + 1.632800102234e-01*V(u2c_17)
+ + -7.710485160351e-02*V(u2c_18) + 1.817059814930e-01*V(u2c_19))
B_u3_15 u3_15 0 V = tanh_psi(0.0 + 2.046545445919e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.561491489410e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.512126624584e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -9.328781068325e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -6.629116833210e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.918087154627e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 1.690723299980e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.809618473053e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 1.717540323734e-01*(V(u2a_8) + (-1)*V(u2b_8)) + -1.412975490093e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.557241529226e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 2.436295151711e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 3.223964571953e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -1.292686164379e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + -1.195086389780e-01*(V(u2a_14) + (-1)*V(u2b_14)) + -1.233121305704e-01*(V(u2a_15) + (-1)*V(u2b_15))
+ + -2.078325748444e-01*(V(u2a_16) + (-1)*V(u2b_16)) + -2.036947906017e-01*(V(u2a_17) + (-1)*V(u2b_17))
+ + -2.057400494814e-01*(V(u2a_18) + (-1)*V(u2b_18)) + 6.975707411766e-02*(V(u2a_19) + (-1)*V(u2b_19)) + 2.620597183704e-02*V(u2c_0)
+ + -1.799465715885e-01*V(u2c_1) + 1.857315599918e-01*V(u2c_2) + 5.296802520752e-02*V(u2c_3) + -8.520731329918e-02*V(u2c_4)
+ + 1.323379278183e-01*V(u2c_5) + 7.859432697296e-02*V(u2c_6) + -1.599882543087e-02*V(u2c_7) + -4.084362089634e-02*V(u2c_8)
+ + 1.736423075199e-01*V(u2c_9) + -2.062013745308e-01*V(u2c_10) + 2.051138579845e-01*V(u2c_11) + -1.183913201094e-01*V(u2c_12)
+ + -8.933404088020e-02*V(u2c_13) + -2.131734788418e-02*V(u2c_14) + 3.181511163712e-02*V(u2c_15) + -4.055775702000e-02*V(u2c_16)
+ + -8.871452510357e-02*V(u2c_17) + -2.178249806166e-01*V(u2c_18) + -1.662779301405e-01*V(u2c_19))
B_u3_16 u3_16 0 V = tanh_psi(0.0 + -1.120167002082e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 8.710089325905e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + 3.916347026825e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 1.170660257339e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 9.739565849304e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 1.595195531845e-01*(V(u2a_5) + (-1)*V(u2b_5)) + -9.649029374123e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 4.614028334618e-02*(V(u2a_7) + (-1)*V(u2b_7)) + -2.109823524952e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.393219232559e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 9.123265743256e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.806767284870e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 2.561031281948e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 1.221857666969e-01*(V(u2a_13) + (-1)*V(u2b_13)) + -5.409538745880e-03*(V(u2a_14)
+ + (-1)*V(u2b_14)) + 7.122910022736e-02*(V(u2a_15) + (-1)*V(u2b_15)) + -1.111755967140e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + 4.181402921677e-02*(V(u2a_17) + (-1)*V(u2b_17)) + -5.121847987175e-02*(V(u2a_18) + (-1)*V(u2b_18)) + 1.379444897175e-01*(V(u2a_19)
+ + (-1)*V(u2b_19)) + -1.557469218969e-01*V(u2c_0) + 1.916261911392e-01*V(u2c_1) + -1.244411990047e-01*V(u2c_2)
+ + 2.132099568844e-01*V(u2c_3) + -2.141622304916e-01*V(u2c_4) + 6.516414880753e-02*V(u2c_5) + -9.503298997879e-02*V(u2c_6)
+ + 1.651583313942e-01*V(u2c_7) + 6.095603108406e-02*V(u2c_8) + -1.972968876362e-01*V(u2c_9) + 5.897012352943e-02*V(u2c_10)
+ + 1.877400279045e-01*V(u2c_11) + 5.829417705536e-02*V(u2c_12) + -8.851620554924e-02*V(u2c_13) + -1.219639182091e-01*V(u2c_14)
+ + -2.123857289553e-01*V(u2c_15) + -1.469102352858e-01*V(u2c_16) + 1.886373758316e-01*V(u2c_17) + 1.008625328541e-02*V(u2c_18)
+ + 1.282844543457e-01*V(u2c_19))
B_u3_17 u3_17 0 V = tanh_psi(0.0 + 9.210494160652e-02*(V(u2a_0) + (-1)*V(u2b_0)) + 2.116010785103e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 2.118497192860e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -1.677897274494e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 1.557265818119e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 1.178412735462e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 7.689172029495e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.247715726495e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -1.288906931877e-01*(V(u2a_8) + (-1)*V(u2b_8)) + -1.635160744190e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 1.008209586143e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -2.229749113321e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.509724259377e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 1.647270321846e-01*(V(u2a_13) + (-1)*V(u2b_13)) + 9.894427657127e-02*(V(u2a_14)
+ + (-1)*V(u2b_14)) + 1.802507340908e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 1.030125021935e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + -2.074207365513e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -2.063322961330e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + -8.704012632370e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -2.215749472380e-01*V(u2c_0) + 5.929163098335e-02*V(u2c_1)
+ + -1.378169059753e-01*V(u2c_2) + -3.360895812511e-02*V(u2c_3) + 1.491403281689e-01*V(u2c_4) + 1.779617071152e-01*V(u2c_5)
+ + 1.242750883102e-01*V(u2c_6) + 7.014378905296e-02*V(u2c_7) + 2.155421674252e-01*V(u2c_8) + 1.903116703033e-01*V(u2c_9)
+ + -2.622140944004e-02*V(u2c_10) + 6.601065397263e-02*V(u2c_11) + 4.251161217690e-02*V(u2c_12) + 8.025687932968e-02*V(u2c_13)
+ + -5.442951619625e-02*V(u2c_14) + 5.091536045074e-02*V(u2c_15) + 7.176691293716e-02*V(u2c_16) + -7.463586330414e-02*V(u2c_17)
+ + 5.067172646523e-02*V(u2c_18) + -7.878126204014e-02*V(u2c_19))
B_u3_18 u3_18 0 V = tanh_psi(0.0 + 6.510809063911e-03*(V(u2a_0) + (-1)*V(u2b_0)) + -1.700387746096e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -3.418195247650e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 1.775739789009e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 5.723524093628e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -8.028933405876e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 2.130266427994e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.893820762634e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 9.131717681885e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -1.709802746773e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -7.406456768513e-02*(V(u2a_10) + (-1)*V(u2b_10)) + -2.011827975512e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 7.823744416237e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 8.072733879089e-02*(V(u2a_13) + (-1)*V(u2b_13)) + 2.217629551888e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + 1.828834414482e-01*(V(u2a_15) + (-1)*V(u2b_15)) + -7.793773710728e-02*(V(u2a_16) + (-1)*V(u2b_16))
+ + 4.063060879707e-02*(V(u2a_17) + (-1)*V(u2b_17)) + -1.359311044216e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + -1.739088892937e-01*(V(u2a_19) + (-1)*V(u2b_19)) + -7.639057934284e-02*V(u2c_0) + -5.543574690819e-02*V(u2c_1)
+ + 9.260249137878e-02*V(u2c_2) + -1.512954980135e-01*V(u2c_3) + -1.398552954197e-02*V(u2c_4) + 7.709822058678e-02*V(u2c_5)
+ + 4.505127668381e-03*V(u2c_6) + 1.936453580856e-01*V(u2c_7) + -1.523673087358e-01*V(u2c_8) + 1.718547046185e-01*V(u2c_9)
+ + 1.278997957706e-01*V(u2c_10) + 1.794300973415e-01*V(u2c_11) + -2.161579132080e-01*V(u2c_12) + -1.655716896057e-01*V(u2c_13)
+ + 1.442505717278e-01*V(u2c_14) + 9.534931182861e-02*V(u2c_15) + -5.110616981983e-02*V(u2c_16) + 6.070452928543e-02*V(u2c_17)
+ + -1.515493094921e-01*V(u2c_18) + 4.120132327080e-02*V(u2c_19))
B_u3_19 u3_19 0 V = tanh_psi(0.0 + 1.208142638206e-01*(V(u2a_0) + (-1)*V(u2b_0)) + 6.128406524658e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.612686216831e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 7.324844598770e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -1.156323477626e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -2.678592503071e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 2.164644002914e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 6.136545538902e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 1.279725432396e-01*(V(u2a_8) + (-1)*V(u2b_8)) + -7.517759501934e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 1.195079982281e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 1.191225051880e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 1.630593836308e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -8.957101404667e-02*(V(u2a_13) + (-1)*V(u2b_13)) + 5.001348257065e-02*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -6.756052374840e-02*(V(u2a_15) + (-1)*V(u2b_15)) + -9.458401799202e-02*(V(u2a_16) + (-1)*V(u2b_16))
+ + 1.894714236259e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -2.029668688774e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + -7.436171174049e-03*(V(u2a_19) + (-1)*V(u2b_19)) + 3.485074639320e-02*V(u2c_0) + 1.264717876911e-01*V(u2c_1)
+ + -1.006249859929e-01*V(u2c_2) + 2.007146179676e-02*V(u2c_3) + 6.909495592117e-02*V(u2c_4) + 1.944779157639e-01*V(u2c_5)
+ + 1.814183890820e-01*V(u2c_6) + 1.028218269348e-01*V(u2c_7) + -1.391186714172e-01*V(u2c_8) + -7.676677405834e-02*V(u2c_9)
+ + 2.073499560356e-02*V(u2c_10) + 3.792047500610e-04*V(u2c_11) + -1.758575141430e-01*V(u2c_12) + -1.389964967966e-01*V(u2c_13)
+ + 1.786003112793e-01*V(u2c_14) + -1.338911354542e-01*V(u2c_15) + -1.314748823643e-02*V(u2c_16) + -1.600676476955e-01*V(u2c_17)
+ + 2.011645138264e-01*V(u2c_18) + -1.622833162546e-01*V(u2c_19))
B_u3_20 u3_20 0 V = tanh_psi(0.0 + 3.556746244431e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -1.896195560694e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -4.252459108829e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -1.382486522198e-02*(V(u2a_3) + (-1)*V(u2b_3)) + 1.721191108227e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 9.782859683037e-02*(V(u2a_5) + (-1)*V(u2b_5)) + -1.684455722570e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.118039488792e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 3.319320082664e-02*(V(u2a_8) + (-1)*V(u2b_8)) + 1.011232435703e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.004281863570e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -1.854413747787e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.645573675632e-01*(V(u2a_12) + (-1)*V(u2b_12)) + -2.004885524511e-01*(V(u2a_13) + (-1)*V(u2b_13))
+ + -2.703942358494e-02*(V(u2a_14) + (-1)*V(u2b_14)) + -1.892590671778e-01*(V(u2a_15) + (-1)*V(u2b_15))
+ + -2.048249989748e-01*(V(u2a_16) + (-1)*V(u2b_16)) + -1.271983981133e-02*(V(u2a_17) + (-1)*V(u2b_17))
+ + 3.177314996719e-03*(V(u2a_18) + (-1)*V(u2b_18)) + 1.523025333881e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -7.470415532589e-02*V(u2c_0)
+ + 4.071041941643e-03*V(u2c_1) + 1.544950902462e-01*V(u2c_2) + 1.968041360378e-01*V(u2c_3) + 1.229254007339e-01*V(u2c_4)
+ + 3.532227873802e-02*V(u2c_5) + -1.890589892864e-01*V(u2c_6) + -4.671198129654e-02*V(u2c_7) + -1.805671006441e-01*V(u2c_8)
+ + 1.062788963318e-01*V(u2c_9) + -1.516242921352e-01*V(u2c_10) + 6.854417920113e-02*V(u2c_11) + -2.224648445845e-01*V(u2c_12)
+ + 2.483031153679e-02*V(u2c_13) + -5.008837580681e-02*V(u2c_14) + 6.260904669762e-02*V(u2c_15) + 1.568424701691e-01*V(u2c_16)
+ + -6.308063864708e-02*V(u2c_17) + 1.666752696037e-01*V(u2c_18) + -1.369825303555e-01*V(u2c_19))
B_u3_21 u3_21 0 V = tanh_psi(0.0 + -4.358957707882e-02*(V(u2a_0) + (-1)*V(u2b_0)) + 9.692725539207e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + -2.035661041737e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -1.056314408779e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -1.047748476267e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 2.218003571033e-01*(V(u2a_5) + (-1)*V(u2b_5)) + -1.178903877735e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.466533243656e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 6.123068928719e-02*(V(u2a_8) + (-1)*V(u2b_8)) + 1.258564293385e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 1.131716668606e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -1.032446324825e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + -2.189271450043e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 6.517040729523e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + -2.154197692871e-01*(V(u2a_14) + (-1)*V(u2b_14)) + 2.233469188213e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 7.725977897644e-02*(V(u2a_16)
+ + (-1)*V(u2b_16)) + 1.955811083317e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 1.934709548950e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + -2.208375632763e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 1.698568761349e-01*V(u2c_0) + 1.603538393974e-01*V(u2c_1)
+ + -4.653832316399e-02*V(u2c_2) + -6.126525998116e-02*V(u2c_3) + -1.491235196590e-01*V(u2c_4) + -5.921466648579e-02*V(u2c_5)
+ + 1.986499726772e-01*V(u2c_6) + -1.757080554962e-01*V(u2c_7) + -3.985558450222e-02*V(u2c_8) + -1.797777414322e-01*V(u2c_9)
+ + 1.504312157631e-01*V(u2c_10) + 5.280235409737e-02*V(u2c_11) + -1.791547834873e-01*V(u2c_12) + 1.988320052624e-01*V(u2c_13)
+ + 1.575680971146e-01*V(u2c_14) + -1.232342422009e-01*V(u2c_15) + -3.724944591522e-02*V(u2c_16) + 1.163634657860e-01*V(u2c_17)
+ + -4.929973185062e-02*V(u2c_18) + -2.038887143135e-01*V(u2c_19))
B_u3_22 u3_22 0 V = tanh_psi(0.0 + 5.111080408096e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -4.242503643036e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.199907660484e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 3.803363442421e-02*(V(u2a_3) + (-1)*V(u2b_3)) + 1.069103181362e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -6.937970221043e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 3.335392475128e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.057508587837e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -1.061364933848e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 2.370265126228e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 8.102360367775e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.533071696758e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 1.485716700554e-01*(V(u2a_12) + (-1)*V(u2b_12)) + -7.354269921780e-02*(V(u2a_13) + (-1)*V(u2b_13)) + 1.845584511757e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.617380380630e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 8.962887525558e-02*(V(u2a_16) + (-1)*V(u2b_16))
+ + 1.685262024403e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -3.537204861641e-02*(V(u2a_18) + (-1)*V(u2b_18))
+ + -1.263603270054e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 3.037321567535e-02*V(u2c_0) + -1.958968937397e-01*V(u2c_1)
+ + 6.993269920349e-02*V(u2c_2) + 8.054420351982e-02*V(u2c_3) + -2.788510918617e-02*V(u2c_4) + -1.411363631487e-01*V(u2c_5)
+ + -1.542427986860e-01*V(u2c_6) + -1.113030090928e-01*V(u2c_7) + 2.143714427948e-01*V(u2c_8) + 9.396976232529e-02*V(u2c_9)
+ + -1.336327791214e-01*V(u2c_10) + -6.152443587780e-02*V(u2c_11) + -1.128640398383e-01*V(u2c_12) + -3.218944370747e-02*V(u2c_13)
+ + 1.594442129135e-01*V(u2c_14) + 1.043395698071e-02*V(u2c_15) + 7.712441682816e-02*V(u2c_16) + 1.651904284954e-01*V(u2c_17)
+ + 2.148229479790e-01*V(u2c_18) + 1.115128099918e-01*V(u2c_19))
B_u3_23 u3_23 0 V = tanh_psi(0.0 + 1.819432675838e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -2.102553546429e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 4.424908757210e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -1.059652492404e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 1.609378755093e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 1.230834424496e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 3.898322582245e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.012480258942e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 1.960834264755e-01*(V(u2a_8) + (-1)*V(u2b_8)) + -2.160527706146e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.076053455472e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 2.117113173008e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.364521384239e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 8.143207430840e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + -1.018488183618e-01*(V(u2a_14) + (-1)*V(u2b_14)) + 5.764096975327e-03*(V(u2a_15) + (-1)*V(u2b_15))
+ + -1.950377374887e-01*(V(u2a_16) + (-1)*V(u2b_16)) + -1.303774118423e-01*(V(u2a_17) + (-1)*V(u2b_17))
+ + -1.037769019604e-02*(V(u2a_18) + (-1)*V(u2b_18)) + 1.119548082352e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 5.561658740044e-02*V(u2c_0)
+ + 1.180547773838e-01*V(u2c_1) + -2.968858182430e-02*V(u2c_2) + -2.066486775875e-01*V(u2c_3) + -7.224868237972e-02*V(u2c_4)
+ + -2.612917125225e-02*V(u2c_5) + 2.226704359055e-01*V(u2c_6) + -6.043079495430e-02*V(u2c_7) + 1.114638745785e-01*V(u2c_8)
+ + 7.630294561386e-02*V(u2c_9) + 4.661700129509e-02*V(u2c_10) + -2.168743610382e-01*V(u2c_11) + -1.054824888706e-01*V(u2c_12)
+ + 1.195734739304e-01*V(u2c_13) + 1.726742684841e-01*V(u2c_14) + 6.973010301590e-02*V(u2c_15) + -1.557942330837e-01*V(u2c_16)
+ + 1.363345086575e-01*V(u2c_17) + 2.368003129959e-02*V(u2c_18) + 5.627608299255e-02*V(u2c_19))
B_u3_24 u3_24 0 V = tanh_psi(0.0 + -1.782920658588e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.216943189502e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 2.131584584713e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 1.665180325508e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 8.492982387543e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -5.695383250713e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 8.177569508553e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.666210740805e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -1.198139786720e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.403522193432e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.980957388878e-02*(V(u2a_10) + (-1)*V(u2b_10)) + -1.322817951441e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 1.390529870987e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 1.954803168774e-01*(V(u2a_13) + (-1)*V(u2b_13)) + -6.498718261719e-02*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.084916293621e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 1.947960853577e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + -4.099859297276e-02*(V(u2a_17) + (-1)*V(u2b_17)) + 2.193938791752e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + -1.468929648399e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 8.685711026192e-02*V(u2c_0) + -8.563199639320e-02*V(u2c_1)
+ + -5.410268902779e-03*V(u2c_2) + 8.777916431427e-02*V(u2c_3) + 1.673058569431e-01*V(u2c_4) + 7.075303792953e-02*V(u2c_5)
+ + -4.746067523956e-02*V(u2c_6) + -7.587839663029e-02*V(u2c_7) + -1.945352554321e-02*V(u2c_8) + -1.905107498169e-01*V(u2c_9)
+ + -1.317058205605e-01*V(u2c_10) + 3.402233123779e-03*V(u2c_11) + 2.148972451687e-02*V(u2c_12) + 1.262409985065e-01*V(u2c_13)
+ + -1.649553775787e-01*V(u2c_14) + 2.189755439758e-01*V(u2c_15) + -2.150470167398e-01*V(u2c_16) + -1.586817204952e-01*V(u2c_17)
+ + -4.081578552723e-02*V(u2c_18) + -1.113419011235e-01*V(u2c_19))
B_u3_25 u3_25 0 V = tanh_psi(0.0 + -2.449284493923e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -1.616402417421e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.166933774948e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 1.260510683060e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -8.472460508347e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -2.061321586370e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 1.246678233147e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -5.160875618458e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 3.992798924446e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -1.612222194672e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 2.203749418259e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -2.185660302639e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 3.260329365730e-03*(V(u2a_12) + (-1)*V(u2b_12)) + -1.275906264782e-01*(V(u2a_13) + (-1)*V(u2b_13)) + 1.903145015240e-02*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.352889388800e-01*(V(u2a_15) + (-1)*V(u2b_15)) + -1.859876215458e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + 5.031532049179e-02*(V(u2a_17) + (-1)*V(u2b_17)) + -1.149311587214e-01*(V(u2a_18) + (-1)*V(u2b_18)) + 2.572265267372e-02*(V(u2a_19)
+ + (-1)*V(u2b_19)) + 1.399968266487e-01*V(u2c_0) + 1.169789433479e-01*V(u2c_1) + 1.731906831264e-01*V(u2c_2)
+ + -9.465008974075e-02*V(u2c_3) + 1.532213389874e-01*V(u2c_4) + 1.104451715946e-02*V(u2c_5) + 1.818795502186e-01*V(u2c_6)
+ + -6.915669143200e-02*V(u2c_7) + 2.129039168358e-02*V(u2c_8) + 1.134821176529e-01*V(u2c_9) + -9.095168113708e-02*V(u2c_10)
+ + -1.727645993233e-01*V(u2c_11) + 6.515982747078e-02*V(u2c_12) + -1.357156187296e-01*V(u2c_13) + -1.531690359116e-01*V(u2c_14)
+ + -7.865108549595e-02*V(u2c_15) + 9.920412302017e-02*V(u2c_16) + -2.403298020363e-02*V(u2c_17) + -7.758411765099e-02*V(u2c_18)
+ + -2.167784124613e-01*V(u2c_19))
B_u3_26 u3_26 0 V = tanh_psi(0.0 + -2.129529267550e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.181307360530e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -3.696501255035e-03*(V(u2a_2) + (-1)*V(u2b_2)) + -1.795204728842e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 2.221230268478e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 8.957087993622e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 2.140631973743e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -5.339221656322e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 1.361339390278e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 3.954145312309e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.624404788017e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 4.561436176300e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 9.683695435524e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -1.824807822704e-01*(V(u2a_13) + (-1)*V(u2b_13)) + 1.060024201870e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + 2.006491422653e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 1.399115920067e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + -8.820635080338e-02*(V(u2a_17) + (-1)*V(u2b_17)) + 1.370665132999e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + -1.527370512486e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -1.467972993851e-01*V(u2c_0) + 1.496511697769e-01*V(u2c_1)
+ + 1.179587841034e-01*V(u2c_2) + 2.937865257263e-02*V(u2c_3) + -7.592700421810e-02*V(u2c_4) + 1.911028325558e-01*V(u2c_5)
+ + -2.639530599117e-02*V(u2c_6) + 1.860681176186e-01*V(u2c_7) + 1.627418100834e-01*V(u2c_8) + -2.246201038361e-03*V(u2c_9)
+ + -2.885641157627e-02*V(u2c_10) + -1.968540549278e-01*V(u2c_11) + 1.295645236969e-01*V(u2c_12) + 3.512442111969e-03*V(u2c_13)
+ + 1.622897386551e-02*V(u2c_14) + -1.864954978228e-01*V(u2c_15) + -5.016154050827e-02*V(u2c_16) + -1.806536018848e-01*V(u2c_17)
+ + 2.138752341270e-01*V(u2c_18) + -6.197418272495e-02*V(u2c_19))
B_u3_27 u3_27 0 V = tanh_psi(0.0 + -1.408696919680e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -2.177556157112e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -1.928474903107e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -5.239848792553e-02*(V(u2a_3) + (-1)*V(u2b_3)) + 2.227458953857e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 8.875328302383e-02*(V(u2a_5) + (-1)*V(u2b_5)) + -9.280440211296e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.929163783789e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -2.431817352772e-02*(V(u2a_8) + (-1)*V(u2b_8)) + 4.233226180077e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 5.224663019180e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.252667307854e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -3.301367163658e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -4.315951466560e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + 1.693292260170e-01*(V(u2a_14) + (-1)*V(u2b_14)) + -4.647445678711e-02*(V(u2a_15) + (-1)*V(u2b_15))
+ + -7.436814904213e-02*(V(u2a_16) + (-1)*V(u2b_16)) + -8.855138719082e-02*(V(u2a_17) + (-1)*V(u2b_17))
+ + -1.247091442347e-01*(V(u2a_18) + (-1)*V(u2b_18)) + 2.142976522446e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 2.042904198170e-01*V(u2c_0)
+ + 8.534830808640e-02*V(u2c_1) + -1.156706511974e-01*V(u2c_2) + -1.481697559357e-01*V(u2c_3) + 1.576938927174e-01*V(u2c_4)
+ + 5.166384577751e-02*V(u2c_5) + 4.995948076248e-02*V(u2c_6) + -2.853274345398e-02*V(u2c_7) + 5.624011158943e-03*V(u2c_8)
+ + 1.012158393860e-02*V(u2c_9) + -3.494141995907e-02*V(u2c_10) + -8.570098876953e-02*V(u2c_11) + -1.680068969727e-01*V(u2c_12)
+ + 1.660436391830e-01*V(u2c_13) + -1.155520826578e-01*V(u2c_14) + 3.789201378822e-02*V(u2c_15) + 1.987007558346e-01*V(u2c_16)
+ + 2.733209729195e-02*V(u2c_17) + 9.110307693481e-02*V(u2c_18) + -1.018164306879e-01*V(u2c_19))
B_u3_28 u3_28 0 V = tanh_psi(0.0 + 2.233381569386e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -7.995797693729e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.048799157143e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -7.924811542034e-02*(V(u2a_3) + (-1)*V(u2b_3)) + 4.322832822800e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -3.686077892780e-02*(V(u2a_5) + (-1)*V(u2b_5)) + -1.372398436069e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.028892695904e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -7.750180363655e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -1.704145669937e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -1.628778576851e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -4.520544409752e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 2.157975435257e-01*(V(u2a_12) + (-1)*V(u2b_12)) + -5.875450372696e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + -1.025555729866e-01*(V(u2a_14) + (-1)*V(u2b_14)) + 9.196320176125e-02*(V(u2a_15) + (-1)*V(u2b_15)) + 6.774538755417e-02*(V(u2a_16)
+ + (-1)*V(u2b_16)) + 1.271080672741e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -9.555552899837e-02*(V(u2a_18) + (-1)*V(u2b_18))
+ + 2.120545208454e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 4.410547018051e-02*V(u2c_0) + 1.740114390850e-02*V(u2c_1)
+ + 1.872068345547e-01*V(u2c_2) + 5.398812890053e-02*V(u2c_3) + -1.572603434324e-01*V(u2c_4) + -1.216783300042e-01*V(u2c_5)
+ + -1.310476511717e-01*V(u2c_6) + 9.539619088173e-03*V(u2c_7) + 1.056648194790e-01*V(u2c_8) + 1.969205737114e-01*V(u2c_9)
+ + 2.742946147919e-02*V(u2c_10) + -7.592739164829e-02*V(u2c_11) + -3.023527562618e-02*V(u2c_12) + 1.468865871429e-01*V(u2c_13)
+ + 1.268420815468e-01*V(u2c_14) + -2.156474143267e-01*V(u2c_15) + 1.516659557819e-01*V(u2c_16) + -7.229183614254e-02*V(u2c_17)
+ + -1.463811397552e-01*V(u2c_18) + 1.944455802441e-01*V(u2c_19))
B_u3_29 u3_29 0 V = tanh_psi(0.0 + -1.509177833796e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.871407032013e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + -2.874426543713e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 2.131060361862e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -7.379245758057e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.262162774801e-01*(V(u2a_5) + (-1)*V(u2b_5)) + -1.555427312851e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 8.241063356400e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 2.369101345539e-02*(V(u2a_8) + (-1)*V(u2b_8)) + 1.334477663040e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -9.554091095924e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.435341238976e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.596795618534e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 4.181608557701e-03*(V(u2a_13) + (-1)*V(u2b_13))
+ + -4.451513290405e-02*(V(u2a_14) + (-1)*V(u2b_14)) + -4.817217588425e-02*(V(u2a_15) + (-1)*V(u2b_15))
+ + 1.680509448051e-01*(V(u2a_16) + (-1)*V(u2b_16)) + -1.156578063965e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 1.826936602592e-01*(V(u2a_18)
+ + (-1)*V(u2b_18)) + 6.273552775383e-02*(V(u2a_19) + (-1)*V(u2b_19)) + 4.626438021660e-03*V(u2c_0) + 1.396190226078e-01*V(u2c_1)
+ + -6.511227786541e-02*V(u2c_2) + -5.525885522366e-02*V(u2c_3) + 1.256603896618e-01*V(u2c_4) + 1.852472424507e-01*V(u2c_5)
+ + 1.902021467686e-01*V(u2c_6) + 1.374999582767e-01*V(u2c_7) + 8.281156420708e-02*V(u2c_8) + 1.958404183388e-01*V(u2c_9)
+ + -1.074693202972e-01*V(u2c_10) + -1.893370896578e-01*V(u2c_11) + 3.945454955101e-03*V(u2c_12) + -1.654165089130e-01*V(u2c_13)
+ + -6.175698339939e-02*V(u2c_14) + -1.180967763066e-01*V(u2c_15) + 1.476130783558e-01*V(u2c_16) + -1.499019861221e-01*V(u2c_17)
+ + -2.011016905308e-01*V(u2c_18) + 1.065634489059e-01*V(u2c_19))
B_u3_30 u3_30 0 V = tanh_psi(0.0 + 1.852795481682e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -5.321229994297e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + -7.803490757942e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 5.763056874275e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -1.387553960085e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.748381555080e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 2.139985263348e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.724736690521e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -2.011123299599e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -1.942150890827e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -2.049420773983e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -1.917083263397e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 5.327138304710e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -1.049148738384e-01*(V(u2a_13) + (-1)*V(u2b_13))
+ + -1.380208134651e-02*(V(u2a_14) + (-1)*V(u2b_14)) + 2.162296772003e-01*(V(u2a_15) + (-1)*V(u2b_15))
+ + -6.985801458359e-02*(V(u2a_16) + (-1)*V(u2b_16)) + 1.087197363377e-01*(V(u2a_17) + (-1)*V(u2b_17))
+ + -1.120715588331e-01*(V(u2a_18) + (-1)*V(u2b_18)) + -1.722513884306e-01*(V(u2a_19) + (-1)*V(u2b_19)) + 1.534432172775e-01*V(u2c_0)
+ + -1.945176869631e-01*V(u2c_1) + -3.492845594883e-02*V(u2c_2) + -1.499123424292e-01*V(u2c_3) + -2.973406016827e-02*V(u2c_4)
+ + 1.116541624069e-01*V(u2c_5) + -1.353247165680e-01*V(u2c_6) + -1.099546998739e-01*V(u2c_7) + 1.580359637737e-01*V(u2c_8)
+ + -1.195757836103e-01*V(u2c_9) + 1.930077373981e-01*V(u2c_10) + 1.641291677952e-01*V(u2c_11) + 5.057546496391e-02*V(u2c_12)
+ + 2.524732053280e-02*V(u2c_13) + 1.877368390560e-01*V(u2c_14) + -1.692009270191e-01*V(u2c_15) + 1.311269402504e-01*V(u2c_16)
+ + -1.827155500650e-01*V(u2c_17) + 1.094582676888e-01*V(u2c_18) + -1.965140253305e-01*V(u2c_19))
B_u3_31 u3_31 0 V = tanh_psi(0.0 + -1.575929224491e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.982767134905e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.799577474594e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 1.884216070175e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 2.138352692127e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 3.765821456909e-03*(V(u2a_5) + (-1)*V(u2b_5)) + 2.171638906002e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.021027937531e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -1.468026638031e-02*(V(u2a_8) + (-1)*V(u2b_8)) + 1.372726857662e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 1.328382194042e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 1.002859473228e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -8.173544704914e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -3.487591445446e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + 7.856515049934e-02*(V(u2a_14) + (-1)*V(u2b_14)) + 1.670340299606e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 8.132433891296e-02*(V(u2a_16)
+ + (-1)*V(u2b_16)) + 2.198417484760e-02*(V(u2a_17) + (-1)*V(u2b_17)) + 1.214787662029e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + 2.038524150848e-01*(V(u2a_19) + (-1)*V(u2b_19)) + -2.487465739250e-03*V(u2c_0) + -1.624795347452e-01*V(u2c_1)
+ + 1.276880204678e-01*V(u2c_2) + 1.822946369648e-01*V(u2c_3) + 1.551260054111e-01*V(u2c_4) + -8.455042541027e-02*V(u2c_5)
+ + 1.591913402081e-02*V(u2c_6) + -1.628364026546e-01*V(u2c_7) + -7.061058282852e-02*V(u2c_8) + -9.305609762669e-02*V(u2c_9)
+ + 1.202392280102e-01*V(u2c_10) + 1.249961853027e-01*V(u2c_11) + 2.190364897251e-01*V(u2c_12) + 1.286219358444e-01*V(u2c_13)
+ + -1.037240698934e-01*V(u2c_14) + -1.066920012236e-01*V(u2c_15) + 1.243180334568e-01*V(u2c_16) + -6.890103220940e-03*V(u2c_17)
+ + -1.233018934727e-02*V(u2c_18) + -1.971147954464e-01*V(u2c_19))
B_u3_32 u3_32 0 V = tanh_psi(0.0 + -1.131556034088e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -2.086798250675e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 1.562105715275e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -2.922719717026e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -4.423998296261e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -3.888653218746e-02*(V(u2a_5) + (-1)*V(u2b_5)) + -1.042831763625e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -2.084098607302e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -1.718901097775e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 3.356680274010e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 1.488774120808e-01*(V(u2a_10) + (-1)*V(u2b_10)) + 1.630800366402e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.018957793713e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 1.920667290688e-02*(V(u2a_13) + (-1)*V(u2b_13)) + 1.783576011658e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -8.287440240383e-02*(V(u2a_15) + (-1)*V(u2b_15)) + 8.818116784096e-02*(V(u2a_16) + (-1)*V(u2b_16))
+ + -2.190636545420e-01*(V(u2a_17) + (-1)*V(u2b_17)) + -2.289247512817e-02*(V(u2a_18) + (-1)*V(u2b_18))
+ + -5.357822775841e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -1.958446651697e-01*V(u2c_0) + -2.003894150257e-01*V(u2c_1)
+ + -3.834229707718e-02*V(u2c_2) + -9.530586004257e-02*V(u2c_3) + -1.966781467199e-01*V(u2c_4) + 2.108295261860e-02*V(u2c_5)
+ + -1.659275889397e-01*V(u2c_6) + 1.342316865921e-01*V(u2c_7) + -4.287773370743e-02*V(u2c_8) + -1.381067186594e-01*V(u2c_9)
+ + -1.943667531013e-01*V(u2c_10) + -8.787238597870e-02*V(u2c_11) + -1.754335016012e-01*V(u2c_12) + 1.880543828011e-01*V(u2c_13)
+ + -2.120611220598e-01*V(u2c_14) + 2.024942338467e-01*V(u2c_15) + 1.632215678692e-01*V(u2c_16) + 4.674378037453e-02*V(u2c_17)
+ + -7.560154795647e-02*V(u2c_18) + 1.336522400379e-01*V(u2c_19))
B_u3_33 u3_33 0 V = tanh_psi(0.0 + -1.742032766342e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.279939711094e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 2.154990434647e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -1.517724841833e-01*(V(u2a_3) + (-1)*V(u2b_3)) + -1.754825115204e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 2.167598307133e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 1.847938597202e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -1.971310973167e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 8.109614253044e-02*(V(u2a_8) + (-1)*V(u2b_8)) + 1.138069927692e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -2.224051356316e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -2.129599601030e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 1.766654253006e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 1.790783703327e-01*(V(u2a_13) + (-1)*V(u2b_13)) + -1.338664591312e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + 6.122037768364e-02*(V(u2a_15) + (-1)*V(u2b_15)) + 1.126126945019e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + -1.796744465828e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 1.480237841606e-01*(V(u2a_18) + (-1)*V(u2b_18)) + 1.275647282600e-01*(V(u2a_19)
+ + (-1)*V(u2b_19)) + -4.456314444542e-02*V(u2c_0) + -1.664557009935e-01*V(u2c_1) + -7.855792343616e-02*V(u2c_2)
+ + -1.008651852608e-01*V(u2c_3) + 3.041431307793e-02*V(u2c_4) + -9.737722575665e-02*V(u2c_5) + -9.615935385227e-02*V(u2c_6)
+ + -1.710959821939e-01*V(u2c_7) + -1.890495419502e-02*V(u2c_8) + -2.586629986763e-02*V(u2c_9) + 3.657197952271e-02*V(u2c_10)
+ + 1.767449676991e-01*V(u2c_11) + -4.601132869720e-02*V(u2c_12) + -1.148398369551e-01*V(u2c_13) + -2.831630408764e-02*V(u2c_14)
+ + -1.115114092827e-01*V(u2c_15) + 1.429109573364e-01*V(u2c_16) + 1.911999285221e-01*V(u2c_17) + 2.032250463963e-01*V(u2c_18)
+ + 2.166861295700e-01*V(u2c_19))
B_u3_34 u3_34 0 V = tanh_psi(0.0 + -6.966027617455e-02*(V(u2a_0) + (-1)*V(u2b_0)) + 7.800602912903e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + 3.848668932915e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 1.273595690727e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 1.565283536911e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.819773614407e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 8.381736278534e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 4.280254244804e-02*(V(u2a_7) + (-1)*V(u2b_7)) + -2.131926119328e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.240060627460e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -2.016207277775e-01*(V(u2a_10) + (-1)*V(u2b_10)) + -1.395636498928e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -1.237995326519e-01*(V(u2a_12) + (-1)*V(u2b_12)) + 3.388261795044e-02*(V(u2a_13) + (-1)*V(u2b_13))
+ + -1.520075052977e-01*(V(u2a_14) + (-1)*V(u2b_14)) + -1.939352154732e-01*(V(u2a_15) + (-1)*V(u2b_15))
+ + -5.780954658985e-02*(V(u2a_16) + (-1)*V(u2b_16)) + -4.981531202793e-02*(V(u2a_17) + (-1)*V(u2b_17))
+ + 1.950243711472e-01*(V(u2a_18) + (-1)*V(u2b_18)) + -7.330007851124e-02*(V(u2a_19) + (-1)*V(u2b_19)) + 8.186233043671e-02*V(u2c_0)
+ + -3.725816309452e-02*V(u2c_1) + 5.354151129723e-02*V(u2c_2) + -3.706368803978e-02*V(u2c_3) + 1.113789379597e-01*V(u2c_4)
+ + 1.426152884960e-01*V(u2c_5) + -1.483575701714e-01*V(u2c_6) + 1.720809638500e-01*V(u2c_7) + -4.895263910294e-02*V(u2c_8)
+ + 1.299361884594e-01*V(u2c_9) + 1.737314164639e-01*V(u2c_10) + -2.036798000336e-01*V(u2c_11) + 2.221022844315e-01*V(u2c_12)
+ + 2.062642574310e-02*V(u2c_13) + -2.176259011030e-01*V(u2c_14) + 2.325785160065e-02*V(u2c_15) + 1.788231432438e-01*V(u2c_16)
+ + -4.260595142841e-02*V(u2c_17) + -1.522784084082e-01*V(u2c_18) + 5.863717198372e-02*V(u2c_19))
B_u3_35 u3_35 0 V = tanh_psi(0.0 + -1.356394886971e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.146935224533e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -2.694821357727e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 8.150771260262e-03*(V(u2a_3) + (-1)*V(u2b_3)) + -1.499922573566e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -1.184349879622e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 6.035450100899e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 2.894595265388e-03*(V(u2a_7) + (-1)*V(u2b_7)) + -1.670217514038e-02*(V(u2a_8) + (-1)*V(u2b_8)) + 8.162978291512e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -5.940139293671e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.184010207653e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + 1.057534813881e-01*(V(u2a_12) + (-1)*V(u2b_12)) + -1.563981771469e-01*(V(u2a_13) + (-1)*V(u2b_13)) + 1.921263337135e-02*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -8.769688010216e-02*(V(u2a_15) + (-1)*V(u2b_15)) + -1.098118722439e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + 2.130188345909e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 9.239760041237e-02*(V(u2a_18) + (-1)*V(u2b_18)) + -1.034459397197e-01*(V(u2a_19)
+ + (-1)*V(u2b_19)) + -2.493222057819e-02*V(u2c_0) + -2.094654589891e-01*V(u2c_1) + -7.862202823162e-02*V(u2c_2)
+ + -7.317759096622e-02*V(u2c_3) + -9.098590910435e-02*V(u2c_4) + -7.720243930817e-02*V(u2c_5) + 2.191947400570e-02*V(u2c_6)
+ + -1.401916146278e-02*V(u2c_7) + -4.488106071949e-02*V(u2c_8) + 5.265185236931e-02*V(u2c_9) + -1.219893544912e-01*V(u2c_10)
+ + -1.894190758467e-01*V(u2c_11) + 2.232011854649e-01*V(u2c_12) + 6.985279917717e-02*V(u2c_13) + -2.406549453735e-02*V(u2c_14)
+ + 5.118471384048e-02*V(u2c_15) + -9.369400143623e-02*V(u2c_16) + 4.085642099380e-02*V(u2c_17) + 2.235665023327e-01*V(u2c_18)
+ + -2.084210515022e-01*V(u2c_19))
B_u3_36 u3_36 0 V = tanh_psi(0.0 + -7.235012948513e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -1.286647915840e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -2.042733132839e-02*(V(u2a_2) + (-1)*V(u2b_2)) + 5.283191800117e-02*(V(u2a_3) + (-1)*V(u2b_3)) + 7.190981507301e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 7.171598076820e-02*(V(u2a_5) + (-1)*V(u2b_5)) + -6.898838281631e-02*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.219615936279e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -7.392072677612e-02*(V(u2a_8) + (-1)*V(u2b_8)) + -1.087043136358e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 4.087015986443e-02*(V(u2a_10) + (-1)*V(u2b_10)) + -7.689565420151e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 9.376886487007e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 5.534961819649e-02*(V(u2a_13) + (-1)*V(u2b_13)) + -1.059984415770e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.254007816315e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 2.043795883656e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + -2.847924828529e-03*(V(u2a_17) + (-1)*V(u2b_17)) + -2.041575908661e-01*(V(u2a_18) + (-1)*V(u2b_18))
+ + 4.296544194221e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -1.948143541813e-01*V(u2c_0) + -1.501642763615e-01*V(u2c_1)
+ + 1.031094193459e-01*V(u2c_2) + -1.106659024954e-01*V(u2c_3) + 7.641214132309e-02*V(u2c_4) + 1.425018310547e-01*V(u2c_5)
+ + -7.364884018898e-02*V(u2c_6) + 1.325427889824e-01*V(u2c_7) + -1.419046223164e-01*V(u2c_8) + -1.916711926460e-01*V(u2c_9)
+ + -1.285055875778e-01*V(u2c_10) + -8.688449859619e-03*V(u2c_11) + 6.871551275253e-03*V(u2c_12) + 2.704042196274e-02*V(u2c_13)
+ + -2.049113959074e-01*V(u2c_14) + -8.742928504944e-03*V(u2c_15) + 8.438605070114e-02*V(u2c_16) + -8.436669409275e-02*V(u2c_17)
+ + 7.259908318520e-02*V(u2c_18) + 6.507393717766e-02*V(u2c_19))
B_u3_37 u3_37 0 V = tanh_psi(0.0 + 1.239431798458e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.330018341541e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + 2.051106691360e-01*(V(u2a_2) + (-1)*V(u2b_2)) + -1.036816835403e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -5.061988532543e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + 1.910087764263e-01*(V(u2a_5) + (-1)*V(u2b_5)) + 1.297727525234e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 1.456137001514e-01*(V(u2a_7) + (-1)*V(u2b_7)) + -2.223235964775e-01*(V(u2a_8) + (-1)*V(u2b_8)) + -1.618629544973e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -4.970446228981e-03*(V(u2a_10) + (-1)*V(u2b_10)) + 1.120411753654e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -6.444896757603e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -1.669389009476e-01*(V(u2a_13) + (-1)*V(u2b_13))
+ + -3.247548639774e-02*(V(u2a_14) + (-1)*V(u2b_14)) + 1.608298718929e-02*(V(u2a_15) + (-1)*V(u2b_15)) + 1.506931483746e-01*(V(u2a_16)
+ + (-1)*V(u2b_16)) + 3.747180104256e-02*(V(u2a_17) + (-1)*V(u2b_17)) + -2.523690462112e-03*(V(u2a_18) + (-1)*V(u2b_18))
+ + 3.040540218353e-02*(V(u2a_19) + (-1)*V(u2b_19)) + -1.878868341446e-01*V(u2c_0) + -5.726006627083e-02*V(u2c_1)
+ + -7.226254045963e-02*V(u2c_2) + 2.094525694847e-01*V(u2c_3) + 1.553326845169e-03*V(u2c_4) + 1.022344231606e-01*V(u2c_5)
+ + 1.993993818760e-01*V(u2c_6) + 1.753300726414e-01*V(u2c_7) + -7.382938265800e-02*V(u2c_8) + -1.797077655792e-01*V(u2c_9)
+ + 1.456781625748e-01*V(u2c_10) + -1.565853655338e-01*V(u2c_11) + -8.156879246235e-02*V(u2c_12) + -1.354058086872e-01*V(u2c_13)
+ + -1.210308298469e-01*V(u2c_14) + 1.558375358582e-01*V(u2c_15) + 9.283423423767e-02*V(u2c_16) + -1.412180662155e-01*V(u2c_17)
+ + 1.443906426430e-01*V(u2c_18) + -1.506660133600e-01*V(u2c_19))
B_u3_38 u3_38 0 V = tanh_psi(0.0 + 8.357176184654e-02*(V(u2a_0) + (-1)*V(u2b_0)) + -1.917418539524e-01*(V(u2a_1) + (-1)*V(u2b_1))
+ + -8.928659558296e-02*(V(u2a_2) + (-1)*V(u2b_2)) + -7.804374396801e-02*(V(u2a_3) + (-1)*V(u2b_3)) + -1.456322968006e-01*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -5.568765103817e-02*(V(u2a_5) + (-1)*V(u2b_5)) + -1.513126492500e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + -2.005796879530e-01*(V(u2a_7) + (-1)*V(u2b_7)) + 1.652711331844e-01*(V(u2a_8) + (-1)*V(u2b_8)) + 1.420238018036e-01*(V(u2a_9)
+ + (-1)*V(u2b_9)) + 4.697674512863e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 9.888470172882e-02*(V(u2a_11) + (-1)*V(u2b_11))
+ + 3.573340177536e-02*(V(u2a_12) + (-1)*V(u2b_12)) + -6.744535267353e-02*(V(u2a_13) + (-1)*V(u2b_13)) + 2.145655453205e-01*(V(u2a_14)
+ + (-1)*V(u2b_14)) + -1.069242283702e-01*(V(u2a_15) + (-1)*V(u2b_15)) + 1.945843398571e-01*(V(u2a_16) + (-1)*V(u2b_16))
+ + 1.793076395988e-01*(V(u2a_17) + (-1)*V(u2b_17)) + 1.120518743992e-01*(V(u2a_18) + (-1)*V(u2b_18)) + 1.764589548111e-01*(V(u2a_19)
+ + (-1)*V(u2b_19)) + 1.538040041924e-01*V(u2c_0) + 8.615213632584e-02*V(u2c_1) + -1.848576962948e-01*V(u2c_2)
+ + -2.871087193489e-02*V(u2c_3) + -1.153138875961e-01*V(u2c_4) + 5.445718765259e-02*V(u2c_5) + -3.255452215672e-02*V(u2c_6)
+ + -2.082503288984e-01*V(u2c_7) + 1.647572517395e-01*V(u2c_8) + -6.157566606998e-02*V(u2c_9) + 5.542853474617e-02*V(u2c_10)
+ + 7.155200839043e-02*V(u2c_11) + 1.175327301025e-01*V(u2c_12) + 1.626443862915e-01*V(u2c_13) + 2.200195193291e-01*V(u2c_14)
+ + 2.191025018692e-01*V(u2c_15) + 1.596838533878e-01*V(u2c_16) + -1.360964030027e-01*V(u2c_17) + 1.508084535599e-01*V(u2c_18)
+ + 1.167323887348e-01*V(u2c_19))
B_u3_39 u3_39 0 V = tanh_psi(0.0 + 1.252652704716e-01*(V(u2a_0) + (-1)*V(u2b_0)) + -1.112878322601e-02*(V(u2a_1) + (-1)*V(u2b_1))
+ + -2.184486240149e-01*(V(u2a_2) + (-1)*V(u2b_2)) + 1.593107879162e-01*(V(u2a_3) + (-1)*V(u2b_3)) + 2.501004934311e-02*(V(u2a_4)
+ + (-1)*V(u2b_4)) + -2.040986716747e-02*(V(u2a_5) + (-1)*V(u2b_5)) + 2.038832008839e-01*(V(u2a_6) + (-1)*V(u2b_6))
+ + 8.108782768250e-02*(V(u2a_7) + (-1)*V(u2b_7)) + 1.697699129581e-01*(V(u2a_8) + (-1)*V(u2b_8)) + -7.129369676113e-02*(V(u2a_9)
+ + (-1)*V(u2b_9)) + -7.354211807251e-02*(V(u2a_10) + (-1)*V(u2b_10)) + 1.010904014111e-01*(V(u2a_11) + (-1)*V(u2b_11))
+ + -9.743964672089e-02*(V(u2a_12) + (-1)*V(u2b_12)) + 2.215383052826e-01*(V(u2a_13) + (-1)*V(u2b_13))
+ + -2.096336930990e-01*(V(u2a_14) + (-1)*V(u2b_14)) + -2.195901572704e-01*(V(u2a_15) + (-1)*V(u2b_15))
+ + 4.141619801521e-02*(V(u2a_16) + (-1)*V(u2b_16)) + 7.571128010750e-02*(V(u2a_17) + (-1)*V(u2b_17)) + -1.083611175418e-01*(V(u2a_18)
+ + (-1)*V(u2b_18)) + 1.198031902313e-01*(V(u2a_19) + (-1)*V(u2b_19)) + -1.745878458023e-01*V(u2c_0) + -2.043121159077e-01*V(u2c_1)
+ + -1.301383376122e-01*V(u2c_2) + -9.027022123337e-02*V(u2c_3) + -1.146376803517e-01*V(u2c_4) + -2.230732440948e-01*V(u2c_5)
+ + -1.845831274986e-01*V(u2c_6) + 1.112866401672e-02*V(u2c_7) + 7.471257448196e-02*V(u2c_8) + -7.547685503960e-02*V(u2c_9)
+ + -3.185211122036e-02*V(u2c_10) + -8.109559118748e-02*V(u2c_11) + 1.246722638607e-01*V(u2c_12) + -4.750281572342e-02*V(u2c_13)
+ + -1.649656593800e-01*V(u2c_14) + -7.105979323387e-02*V(u2c_15) + 1.995402574539e-02*V(u2c_16) + -1.527482867241e-01*V(u2c_17)
+ + 1.180552840233e-01*V(u2c_18) + 1.412410140038e-01*V(u2c_19))
B_out_0 out0 0 V = (7.278533279896e-02 + -1.918177306652e-02*V(u3_0) + 1.761576533318e-02*V(u3_1) + 3.272438049316e-02*V(u3_2)
+ + -4.830924421549e-02*V(u3_3) + -1.217743381858e-01*V(u3_4) + 6.450331211090e-02*V(u3_5) + -8.589151501656e-02*V(u3_6)
+ + 1.109621971846e-01*V(u3_7) + 1.671046018600e-02*V(u3_8) + 3.494243323803e-02*V(u3_9) + 4.696428775787e-03*V(u3_10)
+ + 1.282100379467e-02*V(u3_11) + -7.595064491034e-02*V(u3_12) + -4.257548600435e-02*V(u3_13) + 7.468670606613e-02*V(u3_14)
+ + 9.121544659138e-02*V(u3_15) + -1.224982216954e-01*V(u3_16) + -1.034156829119e-01*V(u3_17) + -3.625615686178e-02*V(u3_18)
+ + -1.273764520884e-01*V(u3_19) + 1.537367701530e-03*V(u3_20) + -7.373278588057e-02*V(u3_21) + 1.483245939016e-01*V(u3_22)
+ + 5.158035457134e-02*V(u3_23) + -2.754446864128e-02*V(u3_24) + 5.362032353878e-02*V(u3_25) + 3.989726305008e-02*V(u3_26)
+ + -1.152427941561e-01*V(u3_27) + -1.805098354816e-02*V(u3_28) + 1.197674721479e-01*V(u3_29) + -9.045767784119e-02*V(u3_30)
+ + 1.073677837849e-02*V(u3_31) + 8.694645762444e-02*V(u3_32) + 6.511779129505e-02*V(u3_33) + -7.530947029591e-02*V(u3_34)
+ + -1.100341603160e-01*V(u3_35) + -2.313059568405e-02*V(u3_36) + -3.146025538445e-02*V(u3_37) + 1.569648534060e-01*V(u3_38)
+ + -9.425801038742e-02*V(u3_39))

.ends psi_nn_psinn_burgers
