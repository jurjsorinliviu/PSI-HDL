* ngspice behavioral subcircuit (B-sources)
* Generated from model: PsiNN_laplace
.subckt psi_nn_psinn_laplace in0 in1 out0 vdd vss

* Activation (fallback-friendly): use tanh() if supported by ngspice, else replace with rational approx
.func tanh_psi(x) { tanh(x) }

B_u13_0 u13_0 0 V = tanh_psi(-5.665620565414e-01 + -8.157656192780e-01*V(in0) + 3.668748140335e-01*V(in1))
B_u14_0 u14_0 0 V = tanh_psi(-5.665620565414e-01 + -8.157656192780e-01*V(in0) + (-1)*(3.668748140335e-01*V(in1)))
B_u13_1 u13_1 0 V = tanh_psi(5.053761005402e-01 + -8.688112497330e-01*V(in0) + -6.140457391739e-01*V(in1))
B_u14_1 u14_1 0 V = tanh_psi(5.053761005402e-01 + -8.688112497330e-01*V(in0) + (-1)*(-6.140457391739e-01*V(in1)))
B_u13_2 u13_2 0 V = tanh_psi(-3.724560737610e-01 + 2.057421207428e-02*V(in0) + -4.692682027817e-01*V(in1))
B_u14_2 u14_2 0 V = tanh_psi(-3.724560737610e-01 + 2.057421207428e-02*V(in0) + (-1)*(-4.692682027817e-01*V(in1)))
B_u13_3 u13_3 0 V = tanh_psi(7.214748859406e-01 + 1.038964986801e-01*V(in0) + 4.739869832993e-01*V(in1))
B_u14_3 u14_3 0 V = tanh_psi(7.214748859406e-01 + 1.038964986801e-01*V(in0) + (-1)*(4.739869832993e-01*V(in1)))
B_u13_4 u13_4 0 V = tanh_psi(6.953829526901e-01 + -3.372356891632e-01*V(in0) + 2.286871671677e-01*V(in1))
B_u14_4 u14_4 0 V = tanh_psi(6.953829526901e-01 + -3.372356891632e-01*V(in0) + (-1)*(2.286871671677e-01*V(in1)))
B_u13_5 u13_5 0 V = tanh_psi(1.714925765991e-01 + -1.404547691345e-01*V(in0) + -9.102548360825e-01*V(in1))
B_u14_5 u14_5 0 V = tanh_psi(1.714925765991e-01 + -1.404547691345e-01*V(in0) + (-1)*(-9.102548360825e-01*V(in1)))
B_u13_6 u13_6 0 V = tanh_psi(-1.126444339752e-01 + -7.897905111313e-01*V(in0) + 5.154902935028e-01*V(in1))
B_u14_6 u14_6 0 V = tanh_psi(-1.126444339752e-01 + -7.897905111313e-01*V(in0) + (-1)*(5.154902935028e-01*V(in1)))
B_u13_7 u13_7 0 V = tanh_psi(6.030070781708e-01 + 6.916701793671e-01*V(in0) + -2.668412923813e-01*V(in1))
B_u14_7 u14_7 0 V = tanh_psi(6.030070781708e-01 + 6.916701793671e-01*V(in0) + (-1)*(-2.668412923813e-01*V(in1)))
B_u13_8 u13_8 0 V = tanh_psi(4.298877716064e-01 + -9.640698432922e-01*V(in0) + -7.888885736465e-01*V(in1))
B_u14_8 u14_8 0 V = tanh_psi(4.298877716064e-01 + -9.640698432922e-01*V(in0) + (-1)*(-7.888885736465e-01*V(in1)))
B_u13_9 u13_9 0 V = tanh_psi(3.285226821899e-01 + 6.515524387360e-01*V(in0) + -6.140619516373e-01*V(in1))
B_u14_9 u14_9 0 V = tanh_psi(3.285226821899e-01 + 6.515524387360e-01*V(in0) + (-1)*(-6.140619516373e-01*V(in1)))
B_u13_10 u13_10 0 V = tanh_psi(2.992457151413e-01 + 3.717818260193e-01*V(in0) + -3.624230623245e-01*V(in1))
B_u14_10 u14_10 0 V = tanh_psi(2.992457151413e-01 + 3.717818260193e-01*V(in0) + (-1)*(-3.624230623245e-01*V(in1)))
B_u13_11 u13_11 0 V = tanh_psi(-3.891658782959e-01 + 9.932315349579e-02*V(in0) + -6.571027040482e-01*V(in1))
B_u14_11 u14_11 0 V = tanh_psi(-3.891658782959e-01 + 9.932315349579e-02*V(in0) + (-1)*(-6.571027040482e-01*V(in1)))
B_u13_12 u13_12 0 V = tanh_psi(2.766536474228e-01 + -8.720550537109e-01*V(in0) + 5.552325248718e-01*V(in1))
B_u14_12 u14_12 0 V = tanh_psi(2.766536474228e-01 + -8.720550537109e-01*V(in0) + (-1)*(5.552325248718e-01*V(in1)))
B_u13_13 u13_13 0 V = tanh_psi(1.132245063782e-01 + -9.015836715698e-01*V(in0) + -9.238231182098e-01*V(in1))
B_u14_13 u14_13 0 V = tanh_psi(1.132245063782e-01 + -9.015836715698e-01*V(in0) + (-1)*(-9.238231182098e-01*V(in1)))
B_u13_14 u13_14 0 V = tanh_psi(3.199168443680e-01 + -6.510341167450e-02*V(in0) + -8.745965957642e-01*V(in1))
B_u14_14 u14_14 0 V = tanh_psi(3.199168443680e-01 + -6.510341167450e-02*V(in0) + (-1)*(-8.745965957642e-01*V(in1)))
B_u13_15 u13_15 0 V = tanh_psi(-3.734831809998e-01 + -1.389628648758e-01*V(in0) + -4.848867654800e-01*V(in1))
B_u14_15 u14_15 0 V = tanh_psi(-3.734831809998e-01 + -1.389628648758e-01*V(in0) + (-1)*(-4.848867654800e-01*V(in1)))
B_u13_16 u13_16 0 V = tanh_psi(-2.129594087601e-01 + 7.876802682877e-01*V(in0) + -3.580049276352e-01*V(in1))
B_u14_16 u14_16 0 V = tanh_psi(-2.129594087601e-01 + 7.876802682877e-01*V(in0) + (-1)*(-3.580049276352e-01*V(in1)))
B_u13_17 u13_17 0 V = tanh_psi(-7.329008579254e-01 + -1.050139665604e-01*V(in0) + 4.497967958450e-01*V(in1))
B_u14_17 u14_17 0 V = tanh_psi(-7.329008579254e-01 + -1.050139665604e-01*V(in0) + (-1)*(4.497967958450e-01*V(in1)))
B_u13_18 u13_18 0 V = tanh_psi(8.302590847015e-01 + -8.090028762817e-01*V(in0) + -3.972684144974e-01*V(in1))
B_u14_18 u14_18 0 V = tanh_psi(8.302590847015e-01 + -8.090028762817e-01*V(in0) + (-1)*(-3.972684144974e-01*V(in1)))
B_u13_19 u13_19 0 V = tanh_psi(-6.654369831085e-02 + 7.754015922546e-02*V(in0) + -7.532757520676e-01*V(in1))
B_u14_19 u14_19 0 V = tanh_psi(-6.654369831085e-02 + 7.754015922546e-02*V(in0) + (-1)*(-7.532757520676e-01*V(in1)))
B_u23_0 u23_0 0 V = tanh_psi(-1.732249557972e-01 + -1.069156453013e-01*V(u13_0) + 2.229977846146e-01*V(u13_1) + 1.418948769569e-01*V(u13_2)
+ + 9.682992100716e-02*V(u13_3) + 1.912443637848e-01*V(u13_4) + 1.865863800049e-02*V(u13_5) + 2.017188370228e-01*V(u13_6)
+ + -1.436887979507e-01*V(u13_7) + -1.049832999706e-02*V(u13_8) + -1.834024786949e-01*V(u13_9) + 6.191787123680e-02*V(u13_10)
+ + 1.316170394421e-01*V(u13_11) + 6.485342979431e-02*V(u13_12) + -9.786041080952e-02*V(u13_13) + 1.209068596363e-01*V(u13_14)
+ + 2.027826905251e-01*V(u13_15) + -8.951556682587e-02*V(u13_16) + -1.152959764004e-01*V(u13_17) + -7.188695669174e-02*V(u13_18)
+ + -1.955969780684e-01*V(u13_19) + -1.876783370972e-01*V(u14_0) + -4.335837066174e-02*V(u14_1) + -6.092458963394e-02*V(u14_2)
+ + 1.070877313614e-01*V(u14_3) + 1.768919825554e-02*V(u14_4) + -2.008354961872e-01*V(u14_5) + 2.666249871254e-02*V(u14_6)
+ + 8.711659908295e-02*V(u14_7) + 1.192215681076e-01*V(u14_8) + 2.082380354404e-01*V(u14_9) + 2.548855543137e-02*V(u14_10)
+ + -8.365347981453e-02*V(u14_11) + -5.356708168983e-02*V(u14_12) + 1.709586381912e-01*V(u14_13) + -4.881048202515e-02*V(u14_14)
+ + -9.091950953007e-02*V(u14_15) + -2.043484151363e-01*V(u14_16) + 2.179453969002e-01*V(u14_17) + -5.373707413673e-02*V(u14_18)
+ + 1.592637598515e-02*V(u14_19))
B_u24_0 u24_0 0 V = tanh_psi(-1.732249557972e-01 + -1.876783370972e-01*V(u13_0) + -4.335837066174e-02*V(u13_1) + -6.092458963394e-02*V(u13_2)
+ + 1.070877313614e-01*V(u13_3) + 1.768919825554e-02*V(u13_4) + -2.008354961872e-01*V(u13_5) + 2.666249871254e-02*V(u13_6)
+ + 8.711659908295e-02*V(u13_7) + 1.192215681076e-01*V(u13_8) + 2.082380354404e-01*V(u13_9) + 2.548855543137e-02*V(u13_10)
+ + -8.365347981453e-02*V(u13_11) + -5.356708168983e-02*V(u13_12) + 1.709586381912e-01*V(u13_13) + -4.881048202515e-02*V(u13_14)
+ + -9.091950953007e-02*V(u13_15) + -2.043484151363e-01*V(u13_16) + 2.179453969002e-01*V(u13_17) + -5.373707413673e-02*V(u13_18)
+ + 1.592637598515e-02*V(u13_19) + -1.069156453013e-01*V(u14_0) + 2.229977846146e-01*V(u14_1) + 1.418948769569e-01*V(u14_2)
+ + 9.682992100716e-02*V(u14_3) + 1.912443637848e-01*V(u14_4) + 1.865863800049e-02*V(u14_5) + 2.017188370228e-01*V(u14_6)
+ + -1.436887979507e-01*V(u14_7) + -1.049832999706e-02*V(u14_8) + -1.834024786949e-01*V(u14_9) + 6.191787123680e-02*V(u14_10)
+ + 1.316170394421e-01*V(u14_11) + 6.485342979431e-02*V(u14_12) + -9.786041080952e-02*V(u14_13) + 1.209068596363e-01*V(u14_14)
+ + 2.027826905251e-01*V(u14_15) + -8.951556682587e-02*V(u14_16) + -1.152959764004e-01*V(u14_17) + -7.188695669174e-02*V(u14_18)
+ + -1.955969780684e-01*V(u14_19))
B_u23_1 u23_1 0 V = tanh_psi(-6.416815519333e-02 + -5.015759170055e-02*V(u13_0) + -2.119085192680e-02*V(u13_1) + -2.170503735542e-01*V(u13_2)
+ + 1.008728742599e-01*V(u13_3) + 4.323273897171e-02*V(u13_4) + 1.245056390762e-01*V(u13_5) + 7.585284113884e-02*V(u13_6)
+ + 5.563017725945e-02*V(u13_7) + 9.638354182243e-02*V(u13_8) + 1.615210771561e-01*V(u13_9) + 5.542293190956e-02*V(u13_10)
+ + -2.150042355061e-01*V(u13_11) + -2.607212960720e-02*V(u13_12) + 5.187997221947e-02*V(u13_13) + -6.970798969269e-02*V(u13_14)
+ + 8.932012319565e-02*V(u13_15) + 1.496900320053e-01*V(u13_16) + -2.412851154804e-02*V(u13_17) + 2.432727813721e-02*V(u13_18)
+ + -2.218086570501e-01*V(u13_19) + -1.006783545017e-01*V(u14_0) + -9.573297202587e-02*V(u14_1) + 1.723870635033e-02*V(u14_2)
+ + 1.068624258041e-01*V(u14_3) + 1.110614836216e-01*V(u14_4) + -3.877614438534e-02*V(u14_5) + -1.133689582348e-01*V(u14_6)
+ + -3.567911684513e-02*V(u14_7) + -1.281697750092e-01*V(u14_8) + -1.890425086021e-01*V(u14_9) + 1.145312488079e-01*V(u14_10)
+ + -7.937769591808e-02*V(u14_11) + 2.196837067604e-01*V(u14_12) + -2.523522078991e-02*V(u14_13) + -2.802094817162e-02*V(u14_14)
+ + 3.956255316734e-02*V(u14_15) + -4.957705736160e-02*V(u14_16) + -2.069058120251e-01*V(u14_17) + -9.555327892303e-02*V(u14_18)
+ + -3.399403393269e-02*V(u14_19))
B_u24_1 u24_1 0 V = tanh_psi(-6.416815519333e-02 + -1.006783545017e-01*V(u13_0) + -9.573297202587e-02*V(u13_1) + 1.723870635033e-02*V(u13_2)
+ + 1.068624258041e-01*V(u13_3) + 1.110614836216e-01*V(u13_4) + -3.877614438534e-02*V(u13_5) + -1.133689582348e-01*V(u13_6)
+ + -3.567911684513e-02*V(u13_7) + -1.281697750092e-01*V(u13_8) + -1.890425086021e-01*V(u13_9) + 1.145312488079e-01*V(u13_10)
+ + -7.937769591808e-02*V(u13_11) + 2.196837067604e-01*V(u13_12) + -2.523522078991e-02*V(u13_13) + -2.802094817162e-02*V(u13_14)
+ + 3.956255316734e-02*V(u13_15) + -4.957705736160e-02*V(u13_16) + -2.069058120251e-01*V(u13_17) + -9.555327892303e-02*V(u13_18)
+ + -3.399403393269e-02*V(u13_19) + -5.015759170055e-02*V(u14_0) + -2.119085192680e-02*V(u14_1) + -2.170503735542e-01*V(u14_2)
+ + 1.008728742599e-01*V(u14_3) + 4.323273897171e-02*V(u14_4) + 1.245056390762e-01*V(u14_5) + 7.585284113884e-02*V(u14_6)
+ + 5.563017725945e-02*V(u14_7) + 9.638354182243e-02*V(u14_8) + 1.615210771561e-01*V(u14_9) + 5.542293190956e-02*V(u14_10)
+ + -2.150042355061e-01*V(u14_11) + -2.607212960720e-02*V(u14_12) + 5.187997221947e-02*V(u14_13) + -6.970798969269e-02*V(u14_14)
+ + 8.932012319565e-02*V(u14_15) + 1.496900320053e-01*V(u14_16) + -2.412851154804e-02*V(u14_17) + 2.432727813721e-02*V(u14_18)
+ + -2.218086570501e-01*V(u14_19))
B_u23_2 u23_2 0 V = tanh_psi(-2.753336131573e-01 + 1.895276308060e-01*V(u13_0) + 1.540527045727e-01*V(u13_1) + -1.610676199198e-01*V(u13_2)
+ + -3.934964537621e-03*V(u13_3) + 1.491388678551e-01*V(u13_4) + 1.162090897560e-01*V(u13_5) + -9.158058464527e-02*V(u13_6)
+ + 1.358382701874e-01*V(u13_7) + 3.965309262276e-02*V(u13_8) + -1.837584376335e-01*V(u13_9) + 5.317336320877e-02*V(u13_10)
+ + -6.799779832363e-02*V(u13_11) + 5.633881688118e-02*V(u13_12) + -6.237995624542e-02*V(u13_13) + -2.054966539145e-01*V(u13_14)
+ + -1.630732715130e-01*V(u13_15) + 5.350658297539e-02*V(u13_16) + 1.454523801804e-01*V(u13_17) + -1.373763382435e-02*V(u13_18)
+ + -2.010378986597e-01*V(u13_19) + -2.079397439957e-02*V(u14_0) + 4.638853669167e-02*V(u14_1) + 4.094991087914e-02*V(u14_2)
+ + 2.043009996414e-01*V(u14_3) + 1.345939636230e-01*V(u14_4) + 2.152521312237e-01*V(u14_5) + -2.000673264265e-01*V(u14_6)
+ + -2.142727673054e-01*V(u14_7) + -9.878801554441e-02*V(u14_8) + -1.248012483120e-02*V(u14_9) + 1.323001086712e-01*V(u14_10)
+ + 5.800217390060e-02*V(u14_11) + 1.528589427471e-01*V(u14_12) + -1.836452037096e-01*V(u14_13) + 1.802847981453e-01*V(u14_14)
+ + -2.143193781376e-02*V(u14_15) + 2.650600671768e-02*V(u14_16) + 1.152135133743e-01*V(u14_17) + -5.003687739372e-02*V(u14_18)
+ + -6.913381814957e-02*V(u14_19))
B_u24_2 u24_2 0 V = tanh_psi(-2.753336131573e-01 + -2.079397439957e-02*V(u13_0) + 4.638853669167e-02*V(u13_1) + 4.094991087914e-02*V(u13_2)
+ + 2.043009996414e-01*V(u13_3) + 1.345939636230e-01*V(u13_4) + 2.152521312237e-01*V(u13_5) + -2.000673264265e-01*V(u13_6)
+ + -2.142727673054e-01*V(u13_7) + -9.878801554441e-02*V(u13_8) + -1.248012483120e-02*V(u13_9) + 1.323001086712e-01*V(u13_10)
+ + 5.800217390060e-02*V(u13_11) + 1.528589427471e-01*V(u13_12) + -1.836452037096e-01*V(u13_13) + 1.802847981453e-01*V(u13_14)
+ + -2.143193781376e-02*V(u13_15) + 2.650600671768e-02*V(u13_16) + 1.152135133743e-01*V(u13_17) + -5.003687739372e-02*V(u13_18)
+ + -6.913381814957e-02*V(u13_19) + 1.895276308060e-01*V(u14_0) + 1.540527045727e-01*V(u14_1) + -1.610676199198e-01*V(u14_2)
+ + -3.934964537621e-03*V(u14_3) + 1.491388678551e-01*V(u14_4) + 1.162090897560e-01*V(u14_5) + -9.158058464527e-02*V(u14_6)
+ + 1.358382701874e-01*V(u14_7) + 3.965309262276e-02*V(u14_8) + -1.837584376335e-01*V(u14_9) + 5.317336320877e-02*V(u14_10)
+ + -6.799779832363e-02*V(u14_11) + 5.633881688118e-02*V(u14_12) + -6.237995624542e-02*V(u14_13) + -2.054966539145e-01*V(u14_14)
+ + -1.630732715130e-01*V(u14_15) + 5.350658297539e-02*V(u14_16) + 1.454523801804e-01*V(u14_17) + -1.373763382435e-02*V(u14_18)
+ + -2.010378986597e-01*V(u14_19))
B_u23_3 u23_3 0 V = tanh_psi(-8.109259605408e-02 + -2.956449985504e-02*V(u13_0) + 1.918165087700e-01*V(u13_1) + 2.201344668865e-01*V(u13_2)
+ + 2.507103979588e-02*V(u13_3) + -6.489372253418e-02*V(u13_4) + 4.839172959328e-02*V(u13_5) + -1.542480289936e-01*V(u13_6)
+ + -5.943775177002e-02*V(u13_7) + 1.259253919125e-01*V(u13_8) + 1.167424917221e-01*V(u13_9) + 8.204203844070e-02*V(u13_10)
+ + 1.065957546234e-01*V(u13_11) + -2.324403822422e-02*V(u13_12) + 1.008995473385e-01*V(u13_13) + -6.023791432381e-02*V(u13_14)
+ + 1.015150547028e-01*V(u13_15) + 2.129017412663e-01*V(u13_16) + 8.256429433823e-02*V(u13_17) + -2.310270071030e-02*V(u13_18)
+ + 1.943456828594e-01*V(u13_19) + 1.063197553158e-01*V(u14_0) + 1.767319440842e-02*V(u14_1) + -1.055135652423e-01*V(u14_2)
+ + 1.613362133503e-02*V(u14_3) + 5.276516079903e-02*V(u14_4) + -1.355171650648e-01*V(u14_5) + 1.268017292023e-01*V(u14_6)
+ + 1.370017528534e-01*V(u14_7) + -1.464301049709e-01*V(u14_8) + 6.496301293373e-02*V(u14_9) + 2.027412354946e-01*V(u14_10)
+ + -1.775378286839e-01*V(u14_11) + -1.244495660067e-01*V(u14_12) + -5.932864546776e-02*V(u14_13) + -2.166275680065e-02*V(u14_14)
+ + 9.697633981705e-02*V(u14_15) + 1.495316624641e-03*V(u14_16) + 6.937140226364e-02*V(u14_17) + -2.220125049353e-01*V(u14_18)
+ + -1.754771620035e-01*V(u14_19))
B_u24_3 u24_3 0 V = tanh_psi(-8.109259605408e-02 + 1.063197553158e-01*V(u13_0) + 1.767319440842e-02*V(u13_1) + -1.055135652423e-01*V(u13_2)
+ + 1.613362133503e-02*V(u13_3) + 5.276516079903e-02*V(u13_4) + -1.355171650648e-01*V(u13_5) + 1.268017292023e-01*V(u13_6)
+ + 1.370017528534e-01*V(u13_7) + -1.464301049709e-01*V(u13_8) + 6.496301293373e-02*V(u13_9) + 2.027412354946e-01*V(u13_10)
+ + -1.775378286839e-01*V(u13_11) + -1.244495660067e-01*V(u13_12) + -5.932864546776e-02*V(u13_13) + -2.166275680065e-02*V(u13_14)
+ + 9.697633981705e-02*V(u13_15) + 1.495316624641e-03*V(u13_16) + 6.937140226364e-02*V(u13_17) + -2.220125049353e-01*V(u13_18)
+ + -1.754771620035e-01*V(u13_19) + -2.956449985504e-02*V(u14_0) + 1.918165087700e-01*V(u14_1) + 2.201344668865e-01*V(u14_2)
+ + 2.507103979588e-02*V(u14_3) + -6.489372253418e-02*V(u14_4) + 4.839172959328e-02*V(u14_5) + -1.542480289936e-01*V(u14_6)
+ + -5.943775177002e-02*V(u14_7) + 1.259253919125e-01*V(u14_8) + 1.167424917221e-01*V(u14_9) + 8.204203844070e-02*V(u14_10)
+ + 1.065957546234e-01*V(u14_11) + -2.324403822422e-02*V(u14_12) + 1.008995473385e-01*V(u14_13) + -6.023791432381e-02*V(u14_14)
+ + 1.015150547028e-01*V(u14_15) + 2.129017412663e-01*V(u14_16) + 8.256429433823e-02*V(u14_17) + -2.310270071030e-02*V(u14_18)
+ + 1.943456828594e-01*V(u14_19))
B_u23_4 u23_4 0 V = tanh_psi(-2.924871742725e-01 + -1.168356537819e-01*V(u13_0) + 1.734991669655e-01*V(u13_1) + -6.123261153698e-02*V(u13_2)
+ + -1.082319691777e-01*V(u13_3) + -3.253819048405e-02*V(u13_4) + -1.704099923372e-01*V(u13_5) + 5.691534280777e-02*V(u13_6)
+ + 1.461461186409e-01*V(u13_7) + -1.021445170045e-01*V(u13_8) + -9.253092110157e-02*V(u13_9) + 1.264914870262e-03*V(u13_10)
+ + 1.948104798794e-01*V(u13_11) + 1.648352146149e-01*V(u13_12) + -1.452634632587e-01*V(u13_13) + 1.739301681519e-01*V(u13_14)
+ + -9.757106006145e-02*V(u13_15) + 7.420763373375e-02*V(u13_16) + 1.467452943325e-02*V(u13_17) + -2.137820869684e-01*V(u13_18)
+ + 1.962147355080e-01*V(u13_19) + 2.253068983555e-02*V(u14_0) + 5.332756042480e-02*V(u14_1) + -1.643871217966e-01*V(u14_2)
+ + 2.167261838913e-01*V(u14_3) + -1.691102087498e-01*V(u14_4) + -2.223260998726e-01*V(u14_5) + -1.014180853963e-01*V(u14_6)
+ + -7.980801165104e-02*V(u14_7) + -7.674606144428e-02*V(u14_8) + 1.274342536926e-01*V(u14_9) + 2.042559683323e-01*V(u14_10)
+ + -4.470545053482e-02*V(u14_11) + -9.209935367107e-02*V(u14_12) + 1.690748929977e-01*V(u14_13) + -1.539335846901e-01*V(u14_14)
+ + -9.866635501385e-02*V(u14_15) + -6.075412034988e-03*V(u14_16) + -2.121137678623e-01*V(u14_17) + -6.874054670334e-04*V(u14_18)
+ + 2.043473124504e-01*V(u14_19))
B_u24_4 u24_4 0 V = tanh_psi(-2.924871742725e-01 + 2.253068983555e-02*V(u13_0) + 5.332756042480e-02*V(u13_1) + -1.643871217966e-01*V(u13_2)
+ + 2.167261838913e-01*V(u13_3) + -1.691102087498e-01*V(u13_4) + -2.223260998726e-01*V(u13_5) + -1.014180853963e-01*V(u13_6)
+ + -7.980801165104e-02*V(u13_7) + -7.674606144428e-02*V(u13_8) + 1.274342536926e-01*V(u13_9) + 2.042559683323e-01*V(u13_10)
+ + -4.470545053482e-02*V(u13_11) + -9.209935367107e-02*V(u13_12) + 1.690748929977e-01*V(u13_13) + -1.539335846901e-01*V(u13_14)
+ + -9.866635501385e-02*V(u13_15) + -6.075412034988e-03*V(u13_16) + -2.121137678623e-01*V(u13_17) + -6.874054670334e-04*V(u13_18)
+ + 2.043473124504e-01*V(u13_19) + -1.168356537819e-01*V(u14_0) + 1.734991669655e-01*V(u14_1) + -6.123261153698e-02*V(u14_2)
+ + -1.082319691777e-01*V(u14_3) + -3.253819048405e-02*V(u14_4) + -1.704099923372e-01*V(u14_5) + 5.691534280777e-02*V(u14_6)
+ + 1.461461186409e-01*V(u14_7) + -1.021445170045e-01*V(u14_8) + -9.253092110157e-02*V(u14_9) + 1.264914870262e-03*V(u14_10)
+ + 1.948104798794e-01*V(u14_11) + 1.648352146149e-01*V(u14_12) + -1.452634632587e-01*V(u14_13) + 1.739301681519e-01*V(u14_14)
+ + -9.757106006145e-02*V(u14_15) + 7.420763373375e-02*V(u14_16) + 1.467452943325e-02*V(u14_17) + -2.137820869684e-01*V(u14_18)
+ + 1.962147355080e-01*V(u14_19))
B_u23_5 u23_5 0 V = tanh_psi(-1.296698898077e-01 + 8.350667357445e-02*V(u13_0) + -2.148568034172e-01*V(u13_1) + -1.275949776173e-01*V(u13_2)
+ + -6.329903006554e-02*V(u13_3) + 1.940828263760e-01*V(u13_4) + -7.976447045803e-02*V(u13_5) + -6.765089929104e-02*V(u13_6)
+ + -6.555035710335e-03*V(u13_7) + 1.678435206413e-01*V(u13_8) + -9.147728979588e-02*V(u13_9) + -1.165582984686e-01*V(u13_10)
+ + 9.222733974457e-02*V(u13_11) + -5.669775605202e-02*V(u13_12) + 1.086315512657e-01*V(u13_13) + -2.198500633240e-01*V(u13_14)
+ + 1.478778421879e-01*V(u13_15) + -1.803458780050e-01*V(u13_16) + -1.643686890602e-01*V(u13_17) + -6.734290719032e-02*V(u13_18)
+ + -7.560998201370e-02*V(u13_19) + 1.352894008160e-01*V(u14_0) + -1.392004787922e-01*V(u14_1) + -8.499646186829e-02*V(u14_2)
+ + -8.465023338795e-02*V(u14_3) + 1.241241991520e-01*V(u14_4) + -1.465216279030e-01*V(u14_5) + -1.238263770938e-01*V(u14_6)
+ + -1.422310471535e-01*V(u14_7) + -1.825712919235e-01*V(u14_8) + 1.912286579609e-01*V(u14_9) + -3.373730182648e-02*V(u14_10)
+ + 3.032156825066e-02*V(u14_11) + -2.129949629307e-01*V(u14_12) + -3.218396008015e-02*V(u14_13) + 1.060649752617e-03*V(u14_14)
+ + -1.395415961742e-01*V(u14_15) + 3.876051306725e-02*V(u14_16) + 8.533620834351e-02*V(u14_17) + -4.252354800701e-02*V(u14_18)
+ + -1.828879117966e-01*V(u14_19))
B_u24_5 u24_5 0 V = tanh_psi(-1.296698898077e-01 + 1.352894008160e-01*V(u13_0) + -1.392004787922e-01*V(u13_1) + -8.499646186829e-02*V(u13_2)
+ + -8.465023338795e-02*V(u13_3) + 1.241241991520e-01*V(u13_4) + -1.465216279030e-01*V(u13_5) + -1.238263770938e-01*V(u13_6)
+ + -1.422310471535e-01*V(u13_7) + -1.825712919235e-01*V(u13_8) + 1.912286579609e-01*V(u13_9) + -3.373730182648e-02*V(u13_10)
+ + 3.032156825066e-02*V(u13_11) + -2.129949629307e-01*V(u13_12) + -3.218396008015e-02*V(u13_13) + 1.060649752617e-03*V(u13_14)
+ + -1.395415961742e-01*V(u13_15) + 3.876051306725e-02*V(u13_16) + 8.533620834351e-02*V(u13_17) + -4.252354800701e-02*V(u13_18)
+ + -1.828879117966e-01*V(u13_19) + 8.350667357445e-02*V(u14_0) + -2.148568034172e-01*V(u14_1) + -1.275949776173e-01*V(u14_2)
+ + -6.329903006554e-02*V(u14_3) + 1.940828263760e-01*V(u14_4) + -7.976447045803e-02*V(u14_5) + -6.765089929104e-02*V(u14_6)
+ + -6.555035710335e-03*V(u14_7) + 1.678435206413e-01*V(u14_8) + -9.147728979588e-02*V(u14_9) + -1.165582984686e-01*V(u14_10)
+ + 9.222733974457e-02*V(u14_11) + -5.669775605202e-02*V(u14_12) + 1.086315512657e-01*V(u14_13) + -2.198500633240e-01*V(u14_14)
+ + 1.478778421879e-01*V(u14_15) + -1.803458780050e-01*V(u14_16) + -1.643686890602e-01*V(u14_17) + -6.734290719032e-02*V(u14_18)
+ + -7.560998201370e-02*V(u14_19))
B_u23_6 u23_6 0 V = tanh_psi(1.533342003822e-01 + -2.016437053680e-01*V(u13_0) + 1.316756010056e-03*V(u13_1) + -1.331088840961e-01*V(u13_2)
+ + 6.027758121490e-02*V(u13_3) + 1.342629194260e-01*V(u13_4) + -1.348417103291e-01*V(u13_5) + -1.688975244761e-01*V(u13_6)
+ + 1.366890370846e-01*V(u13_7) + -1.647967696190e-01*V(u13_8) + -6.511113047600e-02*V(u13_9) + 4.442074894905e-02*V(u13_10)
+ + 9.346094727516e-02*V(u13_11) + 8.648264408112e-02*V(u13_12) + 1.216429769993e-01*V(u13_13) + -2.103582024574e-03*V(u13_14)
+ + -5.411404371262e-02*V(u13_15) + 9.234026074409e-02*V(u13_16) + 9.536567330360e-02*V(u13_17) + 8.122521638870e-02*V(u13_18)
+ + 2.918198704720e-02*V(u13_19) + 3.602269291878e-02*V(u14_0) + 1.118198931217e-01*V(u14_1) + 7.519471645355e-02*V(u14_2)
+ + 7.507565617561e-02*V(u14_3) + 1.159795224667e-01*V(u14_4) + 3.984823822975e-02*V(u14_5) + -1.195921748877e-01*V(u14_6)
+ + -7.657900452614e-02*V(u14_7) + 9.657192230225e-02*V(u14_8) + -1.109606400132e-01*V(u14_9) + 7.791200280190e-02*V(u14_10)
+ + 2.002508342266e-01*V(u14_11) + -1.014910936356e-01*V(u14_12) + -2.053037285805e-02*V(u14_13) + -2.991613745689e-02*V(u14_14)
+ + -2.357582747936e-02*V(u14_15) + -9.838767349720e-02*V(u14_16) + -8.065089583397e-03*V(u14_17) + 1.175369620323e-01*V(u14_18)
+ + -1.478721201420e-02*V(u14_19))
B_u24_6 u24_6 0 V = tanh_psi(1.533342003822e-01 + 3.602269291878e-02*V(u13_0) + 1.118198931217e-01*V(u13_1) + 7.519471645355e-02*V(u13_2)
+ + 7.507565617561e-02*V(u13_3) + 1.159795224667e-01*V(u13_4) + 3.984823822975e-02*V(u13_5) + -1.195921748877e-01*V(u13_6)
+ + -7.657900452614e-02*V(u13_7) + 9.657192230225e-02*V(u13_8) + -1.109606400132e-01*V(u13_9) + 7.791200280190e-02*V(u13_10)
+ + 2.002508342266e-01*V(u13_11) + -1.014910936356e-01*V(u13_12) + -2.053037285805e-02*V(u13_13) + -2.991613745689e-02*V(u13_14)
+ + -2.357582747936e-02*V(u13_15) + -9.838767349720e-02*V(u13_16) + -8.065089583397e-03*V(u13_17) + 1.175369620323e-01*V(u13_18)
+ + -1.478721201420e-02*V(u13_19) + -2.016437053680e-01*V(u14_0) + 1.316756010056e-03*V(u14_1) + -1.331088840961e-01*V(u14_2)
+ + 6.027758121490e-02*V(u14_3) + 1.342629194260e-01*V(u14_4) + -1.348417103291e-01*V(u14_5) + -1.688975244761e-01*V(u14_6)
+ + 1.366890370846e-01*V(u14_7) + -1.647967696190e-01*V(u14_8) + -6.511113047600e-02*V(u14_9) + 4.442074894905e-02*V(u14_10)
+ + 9.346094727516e-02*V(u14_11) + 8.648264408112e-02*V(u14_12) + 1.216429769993e-01*V(u14_13) + -2.103582024574e-03*V(u14_14)
+ + -5.411404371262e-02*V(u14_15) + 9.234026074409e-02*V(u14_16) + 9.536567330360e-02*V(u14_17) + 8.122521638870e-02*V(u14_18)
+ + 2.918198704720e-02*V(u14_19))
B_u23_7 u23_7 0 V = tanh_psi(-1.134560853243e-01 + 9.466937184334e-02*V(u13_0) + -2.155687808990e-01*V(u13_1) + -2.602879703045e-02*V(u13_2)
+ + -7.067221403122e-02*V(u13_3) + 2.443313598633e-02*V(u13_4) + 1.289599537849e-01*V(u13_5) + 1.594802737236e-01*V(u13_6)
+ + -8.874726295471e-02*V(u13_7) + -1.049857512116e-01*V(u13_8) + 6.097513437271e-02*V(u13_9) + -1.768895983696e-02*V(u13_10)
+ + 9.418591856956e-02*V(u13_11) + -8.255247771740e-02*V(u13_12) + -1.962505877018e-01*V(u13_13) + 9.520956873894e-02*V(u13_14)
+ + 1.942159831524e-01*V(u13_15) + 1.742480695248e-01*V(u13_16) + -1.130685433745e-01*V(u13_17) + 2.613160014153e-02*V(u13_18)
+ + 1.613665223122e-01*V(u13_19) + 2.905943989754e-02*V(u14_0) + -7.871286571026e-02*V(u14_1) + -3.790068626404e-02*V(u14_2)
+ + 1.728915572166e-01*V(u14_3) + 1.136275529861e-01*V(u14_4) + -1.758023351431e-01*V(u14_5) + 1.805080175400e-01*V(u14_6)
+ + -1.361769288778e-01*V(u14_7) + -7.672332227230e-02*V(u14_8) + 2.090077996254e-01*V(u14_9) + -6.275404989719e-02*V(u14_10)
+ + 4.844218492508e-03*V(u14_11) + -2.936676144600e-02*V(u14_12) + -1.721129417419e-01*V(u14_13) + 1.168784499168e-01*V(u14_14)
+ + 1.667312085629e-01*V(u14_15) + -9.516631066799e-02*V(u14_16) + 9.991341829300e-02*V(u14_17) + 3.752610087395e-02*V(u14_18)
+ + 1.069027185440e-01*V(u14_19))
B_u24_7 u24_7 0 V = tanh_psi(-1.134560853243e-01 + 2.905943989754e-02*V(u13_0) + -7.871286571026e-02*V(u13_1) + -3.790068626404e-02*V(u13_2)
+ + 1.728915572166e-01*V(u13_3) + 1.136275529861e-01*V(u13_4) + -1.758023351431e-01*V(u13_5) + 1.805080175400e-01*V(u13_6)
+ + -1.361769288778e-01*V(u13_7) + -7.672332227230e-02*V(u13_8) + 2.090077996254e-01*V(u13_9) + -6.275404989719e-02*V(u13_10)
+ + 4.844218492508e-03*V(u13_11) + -2.936676144600e-02*V(u13_12) + -1.721129417419e-01*V(u13_13) + 1.168784499168e-01*V(u13_14)
+ + 1.667312085629e-01*V(u13_15) + -9.516631066799e-02*V(u13_16) + 9.991341829300e-02*V(u13_17) + 3.752610087395e-02*V(u13_18)
+ + 1.069027185440e-01*V(u13_19) + 9.466937184334e-02*V(u14_0) + -2.155687808990e-01*V(u14_1) + -2.602879703045e-02*V(u14_2)
+ + -7.067221403122e-02*V(u14_3) + 2.443313598633e-02*V(u14_4) + 1.289599537849e-01*V(u14_5) + 1.594802737236e-01*V(u14_6)
+ + -8.874726295471e-02*V(u14_7) + -1.049857512116e-01*V(u14_8) + 6.097513437271e-02*V(u14_9) + -1.768895983696e-02*V(u14_10)
+ + 9.418591856956e-02*V(u14_11) + -8.255247771740e-02*V(u14_12) + -1.962505877018e-01*V(u14_13) + 9.520956873894e-02*V(u14_14)
+ + 1.942159831524e-01*V(u14_15) + 1.742480695248e-01*V(u14_16) + -1.130685433745e-01*V(u14_17) + 2.613160014153e-02*V(u14_18)
+ + 1.613665223122e-01*V(u14_19))
B_u23_8 u23_8 0 V = tanh_psi(1.091450601816e-01 + 8.160904049873e-02*V(u13_0) + -1.211911663413e-01*V(u13_1) + 2.799332141876e-03*V(u13_2)
+ + -1.014027297497e-01*V(u13_3) + 6.220963597298e-02*V(u13_4) + 4.920169711113e-02*V(u13_5) + -1.530877947807e-01*V(u13_6)
+ + -2.467247843742e-02*V(u13_7) + 3.351792693138e-02*V(u13_8) + -1.252386122942e-01*V(u13_9) + -1.699949502945e-01*V(u13_10)
+ + 1.751749515533e-01*V(u13_11) + 1.945300400257e-01*V(u13_12) + -7.396958768368e-02*V(u13_13) + 1.382251381874e-01*V(u13_14)
+ + 1.298866569996e-01*V(u13_15) + -5.209569633007e-02*V(u13_16) + -1.484320461750e-01*V(u13_17) + 1.980972588062e-01*V(u13_18)
+ + 1.856419742107e-01*V(u13_19) + 1.660691499710e-01*V(u14_0) + -2.052094638348e-01*V(u14_1) + 1.182695627213e-01*V(u14_2)
+ + -7.917627692223e-03*V(u14_3) + -1.802918463945e-01*V(u14_4) + -2.090239524841e-02*V(u14_5) + -9.054531157017e-02*V(u14_6)
+ + -9.121109545231e-02*V(u14_7) + 1.999965906143e-01*V(u14_8) + 1.119387447834e-01*V(u14_9) + -1.599338054657e-01*V(u14_10)
+ + -1.892070025206e-01*V(u14_11) + -1.175957471132e-01*V(u14_12) + -1.646249890327e-01*V(u14_13) + 5.796620249748e-02*V(u14_14)
+ + -1.313091963530e-01*V(u14_15) + 8.364978432655e-02*V(u14_16) + -9.287971258163e-02*V(u14_17) + -1.668457686901e-02*V(u14_18)
+ + 2.708896994591e-03*V(u14_19))
B_u24_8 u24_8 0 V = tanh_psi(1.091450601816e-01 + 1.660691499710e-01*V(u13_0) + -2.052094638348e-01*V(u13_1) + 1.182695627213e-01*V(u13_2)
+ + -7.917627692223e-03*V(u13_3) + -1.802918463945e-01*V(u13_4) + -2.090239524841e-02*V(u13_5) + -9.054531157017e-02*V(u13_6)
+ + -9.121109545231e-02*V(u13_7) + 1.999965906143e-01*V(u13_8) + 1.119387447834e-01*V(u13_9) + -1.599338054657e-01*V(u13_10)
+ + -1.892070025206e-01*V(u13_11) + -1.175957471132e-01*V(u13_12) + -1.646249890327e-01*V(u13_13) + 5.796620249748e-02*V(u13_14)
+ + -1.313091963530e-01*V(u13_15) + 8.364978432655e-02*V(u13_16) + -9.287971258163e-02*V(u13_17) + -1.668457686901e-02*V(u13_18)
+ + 2.708896994591e-03*V(u13_19) + 8.160904049873e-02*V(u14_0) + -1.211911663413e-01*V(u14_1) + 2.799332141876e-03*V(u14_2)
+ + -1.014027297497e-01*V(u14_3) + 6.220963597298e-02*V(u14_4) + 4.920169711113e-02*V(u14_5) + -1.530877947807e-01*V(u14_6)
+ + -2.467247843742e-02*V(u14_7) + 3.351792693138e-02*V(u14_8) + -1.252386122942e-01*V(u14_9) + -1.699949502945e-01*V(u14_10)
+ + 1.751749515533e-01*V(u14_11) + 1.945300400257e-01*V(u14_12) + -7.396958768368e-02*V(u14_13) + 1.382251381874e-01*V(u14_14)
+ + 1.298866569996e-01*V(u14_15) + -5.209569633007e-02*V(u14_16) + -1.484320461750e-01*V(u14_17) + 1.980972588062e-01*V(u14_18)
+ + 1.856419742107e-01*V(u14_19))
B_u23_9 u23_9 0 V = tanh_psi(-1.880507171154e-01 + 6.285506486893e-02*V(u13_0) + -5.013488233089e-02*V(u13_1) + 1.979690194130e-01*V(u13_2)
+ + 2.116891145706e-01*V(u13_3) + -1.698566973209e-01*V(u13_4) + -4.593667387962e-02*V(u13_5) + 1.945950090885e-01*V(u13_6)
+ + 7.288968563080e-02*V(u13_7) + -1.894203126431e-01*V(u13_8) + 9.952735900879e-02*V(u13_9) + 1.090325713158e-01*V(u13_10)
+ + -1.557685732841e-01*V(u13_11) + -4.035501182079e-02*V(u13_12) + -3.131520748138e-02*V(u13_13) + -1.228119432926e-02*V(u13_14)
+ + -2.139724940062e-01*V(u13_15) + -6.247656047344e-02*V(u13_16) + -4.752285778522e-02*V(u13_17) + -8.424529433250e-02*V(u13_18)
+ + 5.506199598312e-02*V(u13_19) + 1.075586080551e-01*V(u14_0) + -1.042935177684e-01*V(u14_1) + 2.009265720844e-01*V(u14_2)
+ + 9.040758013725e-03*V(u14_3) + 9.945827722549e-02*V(u14_4) + -4.074972867966e-02*V(u14_5) + 1.837413907051e-01*V(u14_6)
+ + -5.472150444984e-02*V(u14_7) + 4.069393873215e-02*V(u14_8) + -2.172114104033e-01*V(u14_9) + 5.648216605186e-02*V(u14_10)
+ + 4.000040888786e-02*V(u14_11) + 3.407993912697e-02*V(u14_12) + 1.469527184963e-01*V(u14_13) + -4.380363225937e-02*V(u14_14)
+ + -6.206762790680e-02*V(u14_15) + -1.454943716526e-01*V(u14_16) + -6.314845383167e-02*V(u14_17) + -8.637276291847e-02*V(u14_18)
+ + 2.207036316395e-01*V(u14_19))
B_u24_9 u24_9 0 V = tanh_psi(-1.880507171154e-01 + 1.075586080551e-01*V(u13_0) + -1.042935177684e-01*V(u13_1) + 2.009265720844e-01*V(u13_2)
+ + 9.040758013725e-03*V(u13_3) + 9.945827722549e-02*V(u13_4) + -4.074972867966e-02*V(u13_5) + 1.837413907051e-01*V(u13_6)
+ + -5.472150444984e-02*V(u13_7) + 4.069393873215e-02*V(u13_8) + -2.172114104033e-01*V(u13_9) + 5.648216605186e-02*V(u13_10)
+ + 4.000040888786e-02*V(u13_11) + 3.407993912697e-02*V(u13_12) + 1.469527184963e-01*V(u13_13) + -4.380363225937e-02*V(u13_14)
+ + -6.206762790680e-02*V(u13_15) + -1.454943716526e-01*V(u13_16) + -6.314845383167e-02*V(u13_17) + -8.637276291847e-02*V(u13_18)
+ + 2.207036316395e-01*V(u13_19) + 6.285506486893e-02*V(u14_0) + -5.013488233089e-02*V(u14_1) + 1.979690194130e-01*V(u14_2)
+ + 2.116891145706e-01*V(u14_3) + -1.698566973209e-01*V(u14_4) + -4.593667387962e-02*V(u14_5) + 1.945950090885e-01*V(u14_6)
+ + 7.288968563080e-02*V(u14_7) + -1.894203126431e-01*V(u14_8) + 9.952735900879e-02*V(u14_9) + 1.090325713158e-01*V(u14_10)
+ + -1.557685732841e-01*V(u14_11) + -4.035501182079e-02*V(u14_12) + -3.131520748138e-02*V(u14_13) + -1.228119432926e-02*V(u14_14)
+ + -2.139724940062e-01*V(u14_15) + -6.247656047344e-02*V(u14_16) + -4.752285778522e-02*V(u14_17) + -8.424529433250e-02*V(u14_18)
+ + 5.506199598312e-02*V(u14_19))
B_u23_10 u23_10 0 V = tanh_psi(1.148915588856e-01 + 7.107931375504e-02*V(u13_0) + 3.980055451393e-03*V(u13_1) + 2.765199542046e-02*V(u13_2)
+ + -9.098508954048e-02*V(u13_3) + -6.031492352486e-02*V(u13_4) + 6.316107511520e-02*V(u13_5) + 1.188154816628e-01*V(u13_6)
+ + 3.772228956223e-03*V(u13_7) + -1.799318194389e-02*V(u13_8) + 1.948837339878e-01*V(u13_9) + 1.805701851845e-02*V(u13_10)
+ + -1.678688228130e-01*V(u13_11) + -1.495624780655e-01*V(u13_12) + -2.052568495274e-01*V(u13_13) + 9.738609194756e-03*V(u13_14)
+ + 6.144049763680e-02*V(u13_15) + -6.681488454342e-02*V(u13_16) + 2.016932964325e-01*V(u13_17) + 9.228804707527e-02*V(u13_18)
+ + -1.019677594304e-01*V(u13_19) + 4.161909222603e-02*V(u14_0) + 1.207562386990e-01*V(u14_1) + -1.134648099542e-01*V(u14_2)
+ + -1.508094966412e-01*V(u14_3) + -2.081540375948e-01*V(u14_4) + -1.374473869801e-01*V(u14_5) + -9.572340548038e-02*V(u14_6)
+ + 3.800579905510e-02*V(u14_7) + 1.703767776489e-01*V(u14_8) + -8.378416299820e-03*V(u14_9) + -2.064696997404e-01*V(u14_10)
+ + -1.499106884003e-01*V(u14_11) + 2.085550129414e-01*V(u14_12) + 1.448640525341e-01*V(u14_13) + -1.734601557255e-01*V(u14_14)
+ + -1.415340602398e-01*V(u14_15) + 1.382065713406e-01*V(u14_16) + -6.927984952927e-02*V(u14_17) + 3.320777416229e-02*V(u14_18)
+ + -1.327732503414e-01*V(u14_19))
B_u24_10 u24_10 0 V = tanh_psi(1.148915588856e-01 + 4.161909222603e-02*V(u13_0) + 1.207562386990e-01*V(u13_1) + -1.134648099542e-01*V(u13_2)
+ + -1.508094966412e-01*V(u13_3) + -2.081540375948e-01*V(u13_4) + -1.374473869801e-01*V(u13_5) + -9.572340548038e-02*V(u13_6)
+ + 3.800579905510e-02*V(u13_7) + 1.703767776489e-01*V(u13_8) + -8.378416299820e-03*V(u13_9) + -2.064696997404e-01*V(u13_10)
+ + -1.499106884003e-01*V(u13_11) + 2.085550129414e-01*V(u13_12) + 1.448640525341e-01*V(u13_13) + -1.734601557255e-01*V(u13_14)
+ + -1.415340602398e-01*V(u13_15) + 1.382065713406e-01*V(u13_16) + -6.927984952927e-02*V(u13_17) + 3.320777416229e-02*V(u13_18)
+ + -1.327732503414e-01*V(u13_19) + 7.107931375504e-02*V(u14_0) + 3.980055451393e-03*V(u14_1) + 2.765199542046e-02*V(u14_2)
+ + -9.098508954048e-02*V(u14_3) + -6.031492352486e-02*V(u14_4) + 6.316107511520e-02*V(u14_5) + 1.188154816628e-01*V(u14_6)
+ + 3.772228956223e-03*V(u14_7) + -1.799318194389e-02*V(u14_8) + 1.948837339878e-01*V(u14_9) + 1.805701851845e-02*V(u14_10)
+ + -1.678688228130e-01*V(u14_11) + -1.495624780655e-01*V(u14_12) + -2.052568495274e-01*V(u14_13) + 9.738609194756e-03*V(u14_14)
+ + 6.144049763680e-02*V(u14_15) + -6.681488454342e-02*V(u14_16) + 2.016932964325e-01*V(u14_17) + 9.228804707527e-02*V(u14_18)
+ + -1.019677594304e-01*V(u14_19))
B_u23_11 u23_11 0 V = tanh_psi(3.308436870575e-01 + 4.862123727798e-02*V(u13_0) + 1.059774458408e-01*V(u13_1) + -9.598018229008e-02*V(u13_2)
+ + -1.528137922287e-01*V(u13_3) + 6.681385636330e-02*V(u13_4) + -9.050455689430e-02*V(u13_5) + 5.464354157448e-02*V(u13_6)
+ + -8.941143751144e-03*V(u13_7) + -1.318165659904e-02*V(u13_8) + 5.180579423904e-02*V(u13_9) + 1.403321623802e-01*V(u13_10)
+ + 1.905698180199e-01*V(u13_11) + -1.148592159152e-01*V(u13_12) + 5.734211206436e-02*V(u13_13) + 1.142010986805e-01*V(u13_14)
+ + -1.144297346473e-01*V(u13_15) + -1.476990133524e-01*V(u13_16) + 1.148829162121e-01*V(u13_17) + -5.080930888653e-02*V(u13_18)
+ + 1.532035768032e-01*V(u13_19) + -6.732036173344e-02*V(u14_0) + -6.146553158760e-02*V(u14_1) + -1.714274734259e-01*V(u14_2)
+ + 1.299298107624e-01*V(u14_3) + 5.728077888489e-02*V(u14_4) + 8.737185597420e-02*V(u14_5) + 1.539239287376e-01*V(u14_6)
+ + -1.981125921011e-01*V(u14_7) + 6.648957729340e-02*V(u14_8) + -1.512784361839e-01*V(u14_9) + -4.440821707249e-02*V(u14_10)
+ + -5.509762465954e-02*V(u14_11) + -6.510385870934e-02*V(u14_12) + 1.898910701275e-01*V(u14_13) + -1.449733078480e-01*V(u14_14)
+ + 1.360279917717e-01*V(u14_15) + 2.207593619823e-01*V(u14_16) + -5.201232433319e-02*V(u14_17) + -2.139265835285e-01*V(u14_18)
+ + 4.121392965317e-03*V(u14_19))
B_u24_11 u24_11 0 V = tanh_psi(3.308436870575e-01 + -6.732036173344e-02*V(u13_0) + -6.146553158760e-02*V(u13_1) + -1.714274734259e-01*V(u13_2)
+ + 1.299298107624e-01*V(u13_3) + 5.728077888489e-02*V(u13_4) + 8.737185597420e-02*V(u13_5) + 1.539239287376e-01*V(u13_6)
+ + -1.981125921011e-01*V(u13_7) + 6.648957729340e-02*V(u13_8) + -1.512784361839e-01*V(u13_9) + -4.440821707249e-02*V(u13_10)
+ + -5.509762465954e-02*V(u13_11) + -6.510385870934e-02*V(u13_12) + 1.898910701275e-01*V(u13_13) + -1.449733078480e-01*V(u13_14)
+ + 1.360279917717e-01*V(u13_15) + 2.207593619823e-01*V(u13_16) + -5.201232433319e-02*V(u13_17) + -2.139265835285e-01*V(u13_18)
+ + 4.121392965317e-03*V(u13_19) + 4.862123727798e-02*V(u14_0) + 1.059774458408e-01*V(u14_1) + -9.598018229008e-02*V(u14_2)
+ + -1.528137922287e-01*V(u14_3) + 6.681385636330e-02*V(u14_4) + -9.050455689430e-02*V(u14_5) + 5.464354157448e-02*V(u14_6)
+ + -8.941143751144e-03*V(u14_7) + -1.318165659904e-02*V(u14_8) + 5.180579423904e-02*V(u14_9) + 1.403321623802e-01*V(u14_10)
+ + 1.905698180199e-01*V(u14_11) + -1.148592159152e-01*V(u14_12) + 5.734211206436e-02*V(u14_13) + 1.142010986805e-01*V(u14_14)
+ + -1.144297346473e-01*V(u14_15) + -1.476990133524e-01*V(u14_16) + 1.148829162121e-01*V(u14_17) + -5.080930888653e-02*V(u14_18)
+ + 1.532035768032e-01*V(u14_19))
B_u23_12 u23_12 0 V = tanh_psi(7.031075656414e-02 + -1.852053403854e-02*V(u13_0) + 1.518328487873e-02*V(u13_1) + -8.523394167423e-02*V(u13_2)
+ + 1.080157160759e-01*V(u13_3) + -2.107094973326e-01*V(u13_4) + 4.862534999847e-02*V(u13_5) + -1.300169974566e-01*V(u13_6)
+ + 1.841737627983e-01*V(u13_7) + 1.464917957783e-01*V(u13_8) + -6.291911005974e-03*V(u13_9) + -1.544378697872e-01*V(u13_10)
+ + 1.742309331894e-02*V(u13_11) + 5.018875002861e-03*V(u13_12) + 1.833722889423e-01*V(u13_13) + -1.758245229721e-01*V(u13_14)
+ + -3.342290222645e-02*V(u13_15) + 1.517682075500e-01*V(u13_16) + -1.999523937702e-01*V(u13_17) + 2.142245173454e-01*V(u13_18)
+ + 1.314819455147e-01*V(u13_19) + 4.267182946205e-02*V(u14_0) + 2.868402004242e-02*V(u14_1) + 1.870947480202e-01*V(u14_2)
+ + 2.680298686028e-02*V(u14_3) + -2.227081209421e-01*V(u14_4) + -6.296591460705e-02*V(u14_5) + -8.425627648830e-02*V(u14_6)
+ + -1.180523931980e-01*V(u14_7) + -1.185968667269e-01*V(u14_8) + -1.993906199932e-01*V(u14_9) + 2.981734275818e-02*V(u14_10)
+ + 3.204792737961e-02*V(u14_11) + -1.232761144638e-01*V(u14_12) + -4.274815320969e-02*V(u14_13) + -6.392286717892e-02*V(u14_14)
+ + 4.162442684174e-02*V(u14_15) + -2.641120553017e-02*V(u14_16) + -9.599573910236e-02*V(u14_17) + -1.463704556227e-01*V(u14_18)
+ + -2.129453569651e-01*V(u14_19))
B_u24_12 u24_12 0 V = tanh_psi(7.031075656414e-02 + 4.267182946205e-02*V(u13_0) + 2.868402004242e-02*V(u13_1) + 1.870947480202e-01*V(u13_2)
+ + 2.680298686028e-02*V(u13_3) + -2.227081209421e-01*V(u13_4) + -6.296591460705e-02*V(u13_5) + -8.425627648830e-02*V(u13_6)
+ + -1.180523931980e-01*V(u13_7) + -1.185968667269e-01*V(u13_8) + -1.993906199932e-01*V(u13_9) + 2.981734275818e-02*V(u13_10)
+ + 3.204792737961e-02*V(u13_11) + -1.232761144638e-01*V(u13_12) + -4.274815320969e-02*V(u13_13) + -6.392286717892e-02*V(u13_14)
+ + 4.162442684174e-02*V(u13_15) + -2.641120553017e-02*V(u13_16) + -9.599573910236e-02*V(u13_17) + -1.463704556227e-01*V(u13_18)
+ + -2.129453569651e-01*V(u13_19) + -1.852053403854e-02*V(u14_0) + 1.518328487873e-02*V(u14_1) + -8.523394167423e-02*V(u14_2)
+ + 1.080157160759e-01*V(u14_3) + -2.107094973326e-01*V(u14_4) + 4.862534999847e-02*V(u14_5) + -1.300169974566e-01*V(u14_6)
+ + 1.841737627983e-01*V(u14_7) + 1.464917957783e-01*V(u14_8) + -6.291911005974e-03*V(u14_9) + -1.544378697872e-01*V(u14_10)
+ + 1.742309331894e-02*V(u14_11) + 5.018875002861e-03*V(u14_12) + 1.833722889423e-01*V(u14_13) + -1.758245229721e-01*V(u14_14)
+ + -3.342290222645e-02*V(u14_15) + 1.517682075500e-01*V(u14_16) + -1.999523937702e-01*V(u14_17) + 2.142245173454e-01*V(u14_18)
+ + 1.314819455147e-01*V(u14_19))
B_u23_13 u23_13 0 V = tanh_psi(1.897160708904e-01 + 4.541957378387e-02*V(u13_0) + -3.834132850170e-02*V(u13_1) + 3.204217553139e-02*V(u13_2)
+ + -3.886763751507e-02*V(u13_3) + 3.787943720818e-02*V(u13_4) + 3.897443413734e-02*V(u13_5) + -1.631551831961e-01*V(u13_6)
+ + -1.736758351326e-01*V(u13_7) + 5.595117807388e-03*V(u13_8) + 2.008996903896e-02*V(u13_9) + -8.764541149139e-02*V(u13_10)
+ + -2.114470154047e-01*V(u13_11) + -1.369355022907e-01*V(u13_12) + -4.763439297676e-02*V(u13_13) + -1.473467051983e-01*V(u13_14)
+ + 2.055423259735e-01*V(u13_15) + 6.300085783005e-02*V(u13_16) + -1.023493930697e-01*V(u13_17) + 1.347255706787e-01*V(u13_18)
+ + 1.075607538223e-02*V(u13_19) + -1.332684159279e-01*V(u14_0) + 8.503517508507e-02*V(u14_1) + 1.875781714916e-01*V(u14_2)
+ + 3.818696737289e-02*V(u14_3) + 8.716037869453e-02*V(u14_4) + 1.559898853302e-01*V(u14_5) + 2.116378545761e-01*V(u14_6)
+ + -1.742791384459e-01*V(u14_7) + 1.377215087414e-01*V(u14_8) + 1.735137999058e-01*V(u14_9) + 1.165041327477e-02*V(u14_10)
+ + -2.183405607939e-01*V(u14_11) + 1.887464821339e-01*V(u14_12) + 1.343518197536e-01*V(u14_13) + 1.171556115150e-01*V(u14_14)
+ + 1.874967813492e-01*V(u14_15) + 4.276648163795e-02*V(u14_16) + 1.904137134552e-01*V(u14_17) + -2.014976143837e-01*V(u14_18)
+ + 2.019866406918e-01*V(u14_19))
B_u24_13 u24_13 0 V = tanh_psi(1.897160708904e-01 + -1.332684159279e-01*V(u13_0) + 8.503517508507e-02*V(u13_1) + 1.875781714916e-01*V(u13_2)
+ + 3.818696737289e-02*V(u13_3) + 8.716037869453e-02*V(u13_4) + 1.559898853302e-01*V(u13_5) + 2.116378545761e-01*V(u13_6)
+ + -1.742791384459e-01*V(u13_7) + 1.377215087414e-01*V(u13_8) + 1.735137999058e-01*V(u13_9) + 1.165041327477e-02*V(u13_10)
+ + -2.183405607939e-01*V(u13_11) + 1.887464821339e-01*V(u13_12) + 1.343518197536e-01*V(u13_13) + 1.171556115150e-01*V(u13_14)
+ + 1.874967813492e-01*V(u13_15) + 4.276648163795e-02*V(u13_16) + 1.904137134552e-01*V(u13_17) + -2.014976143837e-01*V(u13_18)
+ + 2.019866406918e-01*V(u13_19) + 4.541957378387e-02*V(u14_0) + -3.834132850170e-02*V(u14_1) + 3.204217553139e-02*V(u14_2)
+ + -3.886763751507e-02*V(u14_3) + 3.787943720818e-02*V(u14_4) + 3.897443413734e-02*V(u14_5) + -1.631551831961e-01*V(u14_6)
+ + -1.736758351326e-01*V(u14_7) + 5.595117807388e-03*V(u14_8) + 2.008996903896e-02*V(u14_9) + -8.764541149139e-02*V(u14_10)
+ + -2.114470154047e-01*V(u14_11) + -1.369355022907e-01*V(u14_12) + -4.763439297676e-02*V(u14_13) + -1.473467051983e-01*V(u14_14)
+ + 2.055423259735e-01*V(u14_15) + 6.300085783005e-02*V(u14_16) + -1.023493930697e-01*V(u14_17) + 1.347255706787e-01*V(u14_18)
+ + 1.075607538223e-02*V(u14_19))
B_u23_14 u23_14 0 V = tanh_psi(-1.554309427738e-01 + -1.833594739437e-01*V(u13_0) + -1.728095412254e-01*V(u13_1) + -1.948737800121e-01*V(u13_2)
+ + 1.091991364956e-01*V(u13_3) + -1.198661327362e-02*V(u13_4) + 8.298826217651e-02*V(u13_5) + 8.483380079269e-03*V(u13_6)
+ + 1.705129444599e-02*V(u13_7) + 8.122655749321e-02*V(u13_8) + -2.107821404934e-02*V(u13_9) + -1.650162786245e-01*V(u13_10)
+ + -4.833798110485e-02*V(u13_11) + -8.786147832870e-02*V(u13_12) + -1.679956912994e-02*V(u13_13) + -1.293655037880e-01*V(u13_14)
+ + -1.609732210636e-01*V(u13_15) + 7.101729512215e-02*V(u13_16) + 1.348165273666e-01*V(u13_17) + -1.699205338955e-01*V(u13_18)
+ + 3.063639998436e-02*V(u13_19) + -2.135698497295e-02*V(u14_0) + -1.850225925446e-01*V(u14_1) + -1.724540293217e-01*V(u14_2)
+ + -1.474786251783e-01*V(u14_3) + 1.992158591747e-02*V(u14_4) + 1.951405107975e-01*V(u14_5) + 1.107752323151e-04*V(u14_6)
+ + 3.477069735527e-02*V(u14_7) + -1.456301361322e-01*V(u14_8) + -7.720139622688e-02*V(u14_9) + -1.343544125557e-01*V(u14_10)
+ + 5.467757582664e-03*V(u14_11) + 5.819925665855e-02*V(u14_12) + 9.716281294823e-02*V(u14_13) + 4.925286769867e-02*V(u14_14)
+ + 9.847253561020e-02*V(u14_15) + -1.277978122234e-01*V(u14_16) + -1.975738704205e-01*V(u14_17) + -1.375943422318e-01*V(u14_18)
+ + 2.205943167210e-01*V(u14_19))
B_u24_14 u24_14 0 V = tanh_psi(-1.554309427738e-01 + -2.135698497295e-02*V(u13_0) + -1.850225925446e-01*V(u13_1) + -1.724540293217e-01*V(u13_2)
+ + -1.474786251783e-01*V(u13_3) + 1.992158591747e-02*V(u13_4) + 1.951405107975e-01*V(u13_5) + 1.107752323151e-04*V(u13_6)
+ + 3.477069735527e-02*V(u13_7) + -1.456301361322e-01*V(u13_8) + -7.720139622688e-02*V(u13_9) + -1.343544125557e-01*V(u13_10)
+ + 5.467757582664e-03*V(u13_11) + 5.819925665855e-02*V(u13_12) + 9.716281294823e-02*V(u13_13) + 4.925286769867e-02*V(u13_14)
+ + 9.847253561020e-02*V(u13_15) + -1.277978122234e-01*V(u13_16) + -1.975738704205e-01*V(u13_17) + -1.375943422318e-01*V(u13_18)
+ + 2.205943167210e-01*V(u13_19) + -1.833594739437e-01*V(u14_0) + -1.728095412254e-01*V(u14_1) + -1.948737800121e-01*V(u14_2)
+ + 1.091991364956e-01*V(u14_3) + -1.198661327362e-02*V(u14_4) + 8.298826217651e-02*V(u14_5) + 8.483380079269e-03*V(u14_6)
+ + 1.705129444599e-02*V(u14_7) + 8.122655749321e-02*V(u14_8) + -2.107821404934e-02*V(u14_9) + -1.650162786245e-01*V(u14_10)
+ + -4.833798110485e-02*V(u14_11) + -8.786147832870e-02*V(u14_12) + -1.679956912994e-02*V(u14_13) + -1.293655037880e-01*V(u14_14)
+ + -1.609732210636e-01*V(u14_15) + 7.101729512215e-02*V(u14_16) + 1.348165273666e-01*V(u14_17) + -1.699205338955e-01*V(u14_18)
+ + 3.063639998436e-02*V(u14_19))
B_u23_15 u23_15 0 V = tanh_psi(-1.266971230507e-02 + 3.580203652382e-02*V(u13_0) + 5.086046457291e-02*V(u13_1) + -6.167800724506e-02*V(u13_2)
+ + -8.590756356716e-02*V(u13_3) + -1.459939926863e-01*V(u13_4) + 1.936781108379e-01*V(u13_5) + 3.414741158485e-02*V(u13_6)
+ + 1.213001012802e-01*V(u13_7) + 1.765666007996e-01*V(u13_8) + -1.986428350210e-01*V(u13_9) + 8.000791072845e-02*V(u13_10)
+ + -1.497850120068e-01*V(u13_11) + -1.786469519138e-01*V(u13_12) + -2.677887678146e-04*V(u13_13) + -3.916209936142e-02*V(u13_14)
+ + 2.727657556534e-03*V(u13_15) + 2.206456065178e-01*V(u13_16) + 5.643132328987e-02*V(u13_17) + 2.752941846848e-02*V(u13_18)
+ + 2.145289480686e-01*V(u13_19) + -1.571333259344e-01*V(u14_0) + -1.989094167948e-01*V(u14_1) + -1.243449673057e-01*V(u14_2)
+ + -2.176359593868e-01*V(u14_3) + 6.079903244972e-02*V(u14_4) + -6.115618348122e-02*V(u14_5) + 1.968171596527e-01*V(u14_6)
+ + -2.016584724188e-01*V(u14_7) + -1.390580683947e-01*V(u14_8) + -6.846392154694e-02*V(u14_9) + -2.047096788883e-01*V(u14_10)
+ + -2.996492385864e-02*V(u14_11) + -1.823681592941e-01*V(u14_12) + -2.219025194645e-01*V(u14_13) + -1.496721804142e-01*V(u14_14)
+ + -1.380860507488e-01*V(u14_15) + 1.269505918026e-01*V(u14_16) + 3.370568156242e-02*V(u14_17) + 6.679981946945e-02*V(u14_18)
+ + 7.226327061653e-02*V(u14_19))
B_u24_15 u24_15 0 V = tanh_psi(-1.266971230507e-02 + -1.571333259344e-01*V(u13_0) + -1.989094167948e-01*V(u13_1) + -1.243449673057e-01*V(u13_2)
+ + -2.176359593868e-01*V(u13_3) + 6.079903244972e-02*V(u13_4) + -6.115618348122e-02*V(u13_5) + 1.968171596527e-01*V(u13_6)
+ + -2.016584724188e-01*V(u13_7) + -1.390580683947e-01*V(u13_8) + -6.846392154694e-02*V(u13_9) + -2.047096788883e-01*V(u13_10)
+ + -2.996492385864e-02*V(u13_11) + -1.823681592941e-01*V(u13_12) + -2.219025194645e-01*V(u13_13) + -1.496721804142e-01*V(u13_14)
+ + -1.380860507488e-01*V(u13_15) + 1.269505918026e-01*V(u13_16) + 3.370568156242e-02*V(u13_17) + 6.679981946945e-02*V(u13_18)
+ + 7.226327061653e-02*V(u13_19) + 3.580203652382e-02*V(u14_0) + 5.086046457291e-02*V(u14_1) + -6.167800724506e-02*V(u14_2)
+ + -8.590756356716e-02*V(u14_3) + -1.459939926863e-01*V(u14_4) + 1.936781108379e-01*V(u14_5) + 3.414741158485e-02*V(u14_6)
+ + 1.213001012802e-01*V(u14_7) + 1.765666007996e-01*V(u14_8) + -1.986428350210e-01*V(u14_9) + 8.000791072845e-02*V(u14_10)
+ + -1.497850120068e-01*V(u14_11) + -1.786469519138e-01*V(u14_12) + -2.677887678146e-04*V(u14_13) + -3.916209936142e-02*V(u14_14)
+ + 2.727657556534e-03*V(u14_15) + 2.206456065178e-01*V(u14_16) + 5.643132328987e-02*V(u14_17) + 2.752941846848e-02*V(u14_18)
+ + 2.145289480686e-01*V(u14_19))
B_u23_16 u23_16 0 V = tanh_psi(-3.037452101707e-01 + 5.365681648254e-02*V(u13_0) + -1.499739289284e-01*V(u13_1) + 1.195328235626e-01*V(u13_2)
+ + 9.889402985573e-02*V(u13_3) + -3.274162113667e-02*V(u13_4) + 1.501476764679e-01*V(u13_5) + 2.241738140583e-02*V(u13_6)
+ + -1.980640441179e-01*V(u13_7) + -4.052011668682e-02*V(u13_8) + 4.526785016060e-02*V(u13_9) + -6.137657165527e-02*V(u13_10)
+ + 1.819289028645e-01*V(u13_11) + 4.951965808868e-02*V(u13_12) + -1.486576497555e-01*V(u13_13) + 1.693002581596e-01*V(u13_14)
+ + -1.750384271145e-01*V(u13_15) + -1.245050951838e-01*V(u13_16) + 2.868872880936e-02*V(u13_17) + 1.596451103687e-01*V(u13_18)
+ + 1.078358888626e-01*V(u13_19) + 2.181246280670e-01*V(u14_0) + -2.036659419537e-01*V(u14_1) + -1.041267588735e-01*V(u14_2)
+ + -1.767677962780e-01*V(u14_3) + 1.667132973671e-02*V(u14_4) + 1.638728380203e-01*V(u14_5) + 3.823354840279e-03*V(u14_6)
+ + -9.344205260277e-03*V(u14_7) + 2.214045822620e-01*V(u14_8) + -1.055996119976e-01*V(u14_9) + -8.238163590431e-02*V(u14_10)
+ + 9.044978022575e-02*V(u14_11) + 1.491578817368e-01*V(u14_12) + -2.052918225527e-01*V(u14_13) + 8.835095167160e-02*V(u14_14)
+ + -1.001143455505e-02*V(u14_15) + -2.081454247236e-01*V(u14_16) + 9.021884202957e-02*V(u14_17) + 1.087427139282e-01*V(u14_18)
+ + 2.180750966072e-01*V(u14_19))
B_u24_16 u24_16 0 V = tanh_psi(-3.037452101707e-01 + 2.181246280670e-01*V(u13_0) + -2.036659419537e-01*V(u13_1) + -1.041267588735e-01*V(u13_2)
+ + -1.767677962780e-01*V(u13_3) + 1.667132973671e-02*V(u13_4) + 1.638728380203e-01*V(u13_5) + 3.823354840279e-03*V(u13_6)
+ + -9.344205260277e-03*V(u13_7) + 2.214045822620e-01*V(u13_8) + -1.055996119976e-01*V(u13_9) + -8.238163590431e-02*V(u13_10)
+ + 9.044978022575e-02*V(u13_11) + 1.491578817368e-01*V(u13_12) + -2.052918225527e-01*V(u13_13) + 8.835095167160e-02*V(u13_14)
+ + -1.001143455505e-02*V(u13_15) + -2.081454247236e-01*V(u13_16) + 9.021884202957e-02*V(u13_17) + 1.087427139282e-01*V(u13_18)
+ + 2.180750966072e-01*V(u13_19) + 5.365681648254e-02*V(u14_0) + -1.499739289284e-01*V(u14_1) + 1.195328235626e-01*V(u14_2)
+ + 9.889402985573e-02*V(u14_3) + -3.274162113667e-02*V(u14_4) + 1.501476764679e-01*V(u14_5) + 2.241738140583e-02*V(u14_6)
+ + -1.980640441179e-01*V(u14_7) + -4.052011668682e-02*V(u14_8) + 4.526785016060e-02*V(u14_9) + -6.137657165527e-02*V(u14_10)
+ + 1.819289028645e-01*V(u14_11) + 4.951965808868e-02*V(u14_12) + -1.486576497555e-01*V(u14_13) + 1.693002581596e-01*V(u14_14)
+ + -1.750384271145e-01*V(u14_15) + -1.245050951838e-01*V(u14_16) + 2.868872880936e-02*V(u14_17) + 1.596451103687e-01*V(u14_18)
+ + 1.078358888626e-01*V(u14_19))
B_u23_17 u23_17 0 V = tanh_psi(1.456266939640e-01 + -7.014682888985e-02*V(u13_0) + -1.405139267445e-01*V(u13_1) + -1.941498070955e-01*V(u13_2)
+ + 5.283981561661e-02*V(u13_3) + 5.949395895004e-02*V(u13_4) + -4.238212108612e-02*V(u13_5) + -1.602634787560e-01*V(u13_6)
+ + 1.056541502476e-01*V(u13_7) + 1.461935043335e-01*V(u13_8) + 2.756637334824e-02*V(u13_9) + -1.751951724291e-01*V(u13_10)
+ + 4.728460311890e-02*V(u13_11) + -6.494656205177e-03*V(u13_12) + -1.298156976700e-01*V(u13_13) + 2.166701257229e-01*V(u13_14)
+ + 3.818047046661e-02*V(u13_15) + 1.303313076496e-01*V(u13_16) + -2.038779407740e-01*V(u13_17) + 1.364978551865e-01*V(u13_18)
+ + 1.029762923717e-01*V(u13_19) + 1.959196925163e-01*V(u14_0) + -1.271742880344e-01*V(u14_1) + -1.484203636646e-01*V(u14_2)
+ + -9.038548171520e-02*V(u14_3) + 1.943687796593e-01*V(u14_4) + 4.251304268837e-02*V(u14_5) + 2.258901298046e-02*V(u14_6)
+ + -1.955258846283e-01*V(u14_7) + 1.368015706539e-01*V(u14_8) + -6.143942475319e-02*V(u14_9) + -1.169224157929e-01*V(u14_10)
+ + -5.089418590069e-02*V(u14_11) + 1.040341258049e-01*V(u14_12) + -5.076470971107e-02*V(u14_13) + 7.964938879013e-02*V(u14_14)
+ + 7.803705334663e-02*V(u14_15) + 8.529803156853e-02*V(u14_16) + 7.822892069817e-02*V(u14_17) + -9.459520876408e-02*V(u14_18)
+ + 5.453312397003e-02*V(u14_19))
B_u24_17 u24_17 0 V = tanh_psi(1.456266939640e-01 + 1.959196925163e-01*V(u13_0) + -1.271742880344e-01*V(u13_1) + -1.484203636646e-01*V(u13_2)
+ + -9.038548171520e-02*V(u13_3) + 1.943687796593e-01*V(u13_4) + 4.251304268837e-02*V(u13_5) + 2.258901298046e-02*V(u13_6)
+ + -1.955258846283e-01*V(u13_7) + 1.368015706539e-01*V(u13_8) + -6.143942475319e-02*V(u13_9) + -1.169224157929e-01*V(u13_10)
+ + -5.089418590069e-02*V(u13_11) + 1.040341258049e-01*V(u13_12) + -5.076470971107e-02*V(u13_13) + 7.964938879013e-02*V(u13_14)
+ + 7.803705334663e-02*V(u13_15) + 8.529803156853e-02*V(u13_16) + 7.822892069817e-02*V(u13_17) + -9.459520876408e-02*V(u13_18)
+ + 5.453312397003e-02*V(u13_19) + -7.014682888985e-02*V(u14_0) + -1.405139267445e-01*V(u14_1) + -1.941498070955e-01*V(u14_2)
+ + 5.283981561661e-02*V(u14_3) + 5.949395895004e-02*V(u14_4) + -4.238212108612e-02*V(u14_5) + -1.602634787560e-01*V(u14_6)
+ + 1.056541502476e-01*V(u14_7) + 1.461935043335e-01*V(u14_8) + 2.756637334824e-02*V(u14_9) + -1.751951724291e-01*V(u14_10)
+ + 4.728460311890e-02*V(u14_11) + -6.494656205177e-03*V(u14_12) + -1.298156976700e-01*V(u14_13) + 2.166701257229e-01*V(u14_14)
+ + 3.818047046661e-02*V(u14_15) + 1.303313076496e-01*V(u14_16) + -2.038779407740e-01*V(u14_17) + 1.364978551865e-01*V(u14_18)
+ + 1.029762923717e-01*V(u14_19))
B_u23_18 u23_18 0 V = tanh_psi(-2.694069147110e-01 + 3.591379523277e-02*V(u13_0) + 5.567058920860e-02*V(u13_1) + -1.967627555132e-01*V(u13_2)
+ + 2.029036879539e-01*V(u13_3) + 1.524528264999e-01*V(u13_4) + -2.123815715313e-01*V(u13_5) + 3.127542138100e-02*V(u13_6)
+ + 1.648958623409e-01*V(u13_7) + -1.867499351501e-01*V(u13_8) + -1.291463077068e-01*V(u13_9) + -3.956812620163e-02*V(u13_10)
+ + 2.163087129593e-01*V(u13_11) + 1.413800120354e-01*V(u13_12) + 1.773874163628e-01*V(u13_13) + -2.064824104309e-01*V(u13_14)
+ + 1.295167207718e-02*V(u13_15) + 9.747147560120e-03*V(u13_16) + 2.003264129162e-01*V(u13_17) + 1.748293638229e-01*V(u13_18)
+ + 3.165638446808e-02*V(u13_19) + 1.513824760914e-01*V(u14_0) + -1.493038386106e-01*V(u14_1) + 1.565249264240e-01*V(u14_2)
+ + -1.313433349133e-01*V(u14_3) + -5.428476631641e-02*V(u14_4) + -1.297919899225e-01*V(u14_5) + -6.986105442047e-02*V(u14_6)
+ + -1.652059406042e-01*V(u14_7) + -1.672624945641e-01*V(u14_8) + -1.121233478189e-01*V(u14_9) + -9.120488166809e-02*V(u14_10)
+ + -1.433756351471e-01*V(u14_11) + -1.605351269245e-01*V(u14_12) + 4.710376262665e-03*V(u14_13) + 2.062373757362e-01*V(u14_14)
+ + 6.226003170013e-04*V(u14_15) + -2.074722051620e-01*V(u14_16) + -1.777251362801e-01*V(u14_17) + -1.852843314409e-01*V(u14_18)
+ + -1.411778628826e-01*V(u14_19))
B_u24_18 u24_18 0 V = tanh_psi(-2.694069147110e-01 + 1.513824760914e-01*V(u13_0) + -1.493038386106e-01*V(u13_1) + 1.565249264240e-01*V(u13_2)
+ + -1.313433349133e-01*V(u13_3) + -5.428476631641e-02*V(u13_4) + -1.297919899225e-01*V(u13_5) + -6.986105442047e-02*V(u13_6)
+ + -1.652059406042e-01*V(u13_7) + -1.672624945641e-01*V(u13_8) + -1.121233478189e-01*V(u13_9) + -9.120488166809e-02*V(u13_10)
+ + -1.433756351471e-01*V(u13_11) + -1.605351269245e-01*V(u13_12) + 4.710376262665e-03*V(u13_13) + 2.062373757362e-01*V(u13_14)
+ + 6.226003170013e-04*V(u13_15) + -2.074722051620e-01*V(u13_16) + -1.777251362801e-01*V(u13_17) + -1.852843314409e-01*V(u13_18)
+ + -1.411778628826e-01*V(u13_19) + 3.591379523277e-02*V(u14_0) + 5.567058920860e-02*V(u14_1) + -1.967627555132e-01*V(u14_2)
+ + 2.029036879539e-01*V(u14_3) + 1.524528264999e-01*V(u14_4) + -2.123815715313e-01*V(u14_5) + 3.127542138100e-02*V(u14_6)
+ + 1.648958623409e-01*V(u14_7) + -1.867499351501e-01*V(u14_8) + -1.291463077068e-01*V(u14_9) + -3.956812620163e-02*V(u14_10)
+ + 2.163087129593e-01*V(u14_11) + 1.413800120354e-01*V(u14_12) + 1.773874163628e-01*V(u14_13) + -2.064824104309e-01*V(u14_14)
+ + 1.295167207718e-02*V(u14_15) + 9.747147560120e-03*V(u14_16) + 2.003264129162e-01*V(u14_17) + 1.748293638229e-01*V(u14_18)
+ + 3.165638446808e-02*V(u14_19))
B_u23_19 u23_19 0 V = tanh_psi(8.421038091183e-02 + -1.222356781363e-01*V(u13_0) + 2.204292118549e-01*V(u13_1) + 9.697338938713e-02*V(u13_2)
+ + 1.527025997639e-01*V(u13_3) + -2.162729501724e-01*V(u13_4) + 1.994348466396e-01*V(u13_5) + -1.138694509864e-01*V(u13_6)
+ + 1.720144152641e-01*V(u13_7) + 6.812605261803e-02*V(u13_8) + 5.991938710213e-02*V(u13_9) + 1.515619754791e-01*V(u13_10)
+ + -1.323441714048e-01*V(u13_11) + -2.533528208733e-02*V(u13_12) + -1.752747297287e-01*V(u13_13) + 2.116901278496e-01*V(u13_14)
+ + -8.060169219971e-02*V(u13_15) + -1.955006271601e-01*V(u13_16) + 1.021742820740e-02*V(u13_17) + -1.522025167942e-01*V(u13_18)
+ + -7.527978718281e-02*V(u13_19) + -8.789032697678e-02*V(u14_0) + -2.705059945583e-02*V(u14_1) + -1.526104658842e-01*V(u14_2)
+ + 1.552372872829e-01*V(u14_3) + 1.705604195595e-01*V(u14_4) + 1.828570663929e-02*V(u14_5) + 1.391230523586e-02*V(u14_6)
+ + 1.303991973400e-01*V(u14_7) + 1.547709107399e-01*V(u14_8) + 8.139789104462e-03*V(u14_9) + -1.058171689510e-02*V(u14_10)
+ + -9.430460631847e-02*V(u14_11) + -8.176109194756e-02*V(u14_12) + -4.337470233440e-02*V(u14_13) + -2.192980051041e-01*V(u14_14)
+ + -4.599955677986e-02*V(u14_15) + 1.484906077385e-01*V(u14_16) + 1.053752005100e-01*V(u14_17) + 2.032355666161e-01*V(u14_18)
+ + 1.680742502213e-01*V(u14_19))
B_u24_19 u24_19 0 V = tanh_psi(8.421038091183e-02 + -8.789032697678e-02*V(u13_0) + -2.705059945583e-02*V(u13_1) + -1.526104658842e-01*V(u13_2)
+ + 1.552372872829e-01*V(u13_3) + 1.705604195595e-01*V(u13_4) + 1.828570663929e-02*V(u13_5) + 1.391230523586e-02*V(u13_6)
+ + 1.303991973400e-01*V(u13_7) + 1.547709107399e-01*V(u13_8) + 8.139789104462e-03*V(u13_9) + -1.058171689510e-02*V(u13_10)
+ + -9.430460631847e-02*V(u13_11) + -8.176109194756e-02*V(u13_12) + -4.337470233440e-02*V(u13_13) + -2.192980051041e-01*V(u13_14)
+ + -4.599955677986e-02*V(u13_15) + 1.484906077385e-01*V(u13_16) + 1.053752005100e-01*V(u13_17) + 2.032355666161e-01*V(u13_18)
+ + 1.680742502213e-01*V(u13_19) + -1.222356781363e-01*V(u14_0) + 2.204292118549e-01*V(u14_1) + 9.697338938713e-02*V(u14_2)
+ + 1.527025997639e-01*V(u14_3) + -2.162729501724e-01*V(u14_4) + 1.994348466396e-01*V(u14_5) + -1.138694509864e-01*V(u14_6)
+ + 1.720144152641e-01*V(u14_7) + 6.812605261803e-02*V(u14_8) + 5.991938710213e-02*V(u14_9) + 1.515619754791e-01*V(u14_10)
+ + -1.323441714048e-01*V(u14_11) + -2.533528208733e-02*V(u14_12) + -1.752747297287e-01*V(u14_13) + 2.116901278496e-01*V(u14_14)
+ + -8.060169219971e-02*V(u14_15) + -1.955006271601e-01*V(u14_16) + 1.021742820740e-02*V(u14_17) + -1.522025167942e-01*V(u14_18)
+ + -7.527978718281e-02*V(u14_19))
B_u32_0 u32_0 0 V = tanh_psi(2.064499258995e-01 + 1.980400681496e-01*(V(u23_0) + V(u24_0)) + -1.081833019853e-01*(V(u23_1) + V(u24_1))
+ + 1.237388551235e-01*(V(u23_2) + V(u24_2)) + -7.644039392471e-02*(V(u23_3) + V(u24_3)) + 2.213596999645e-01*(V(u23_4) + V(u24_4))
+ + 6.528615951538e-03*(V(u23_5) + V(u24_5)) + -2.277734875679e-02*(V(u23_6) + V(u24_6)) + -2.921703457832e-02*(V(u23_7) + V(u24_7))
+ + -6.159272789955e-02*(V(u23_8) + V(u24_8)) + -1.188923493028e-01*(V(u23_9) + V(u24_9)) + -1.992398500443e-02*(V(u23_10)
+ + V(u24_10)) + 8.315867185593e-02*(V(u23_11) + V(u24_11)) + 1.537846028805e-01*(V(u23_12) + V(u24_12))
+ + -1.541674435139e-01*(V(u23_13) + V(u24_13)) + 1.727891266346e-01*(V(u23_14) + V(u24_14)) + -1.922616958618e-01*(V(u23_15)
+ + V(u24_15)) + -1.786346137524e-01*(V(u23_16) + V(u24_16)) + -1.400151252747e-01*(V(u23_17) + V(u24_17))
+ + -9.125387668610e-02*(V(u23_18) + V(u24_18)) + -2.223947942257e-01*(V(u23_19) + V(u24_19)))
B_u32_1 u32_1 0 V = tanh_psi(3.509033918381e-01 + 1.084710061550e-01*(V(u23_0) + V(u24_0)) + 1.708485186100e-02*(V(u23_1) + V(u24_1))
+ + 9.542787075043e-02*(V(u23_2) + V(u24_2)) + -1.652163267136e-01*(V(u23_3) + V(u24_3)) + -2.109819650650e-02*(V(u23_4) + V(u24_4))
+ + -6.784178316593e-02*(V(u23_5) + V(u24_5)) + 6.012013554573e-02*(V(u23_6) + V(u24_6)) + -1.492698043585e-01*(V(u23_7) + V(u24_7))
+ + -2.677793800831e-02*(V(u23_8) + V(u24_8)) + -2.226728498936e-01*(V(u23_9) + V(u24_9)) + -1.249221265316e-01*(V(u23_10)
+ + V(u24_10)) + 3.365239500999e-02*(V(u23_11) + V(u24_11)) + 8.726724982262e-02*(V(u23_12) + V(u24_12))
+ + 1.395924389362e-01*(V(u23_13) + V(u24_13)) + 2.122690081596e-01*(V(u23_14) + V(u24_14)) + 1.578594744205e-02*(V(u23_15)
+ + V(u24_15)) + -9.238401055336e-02*(V(u23_16) + V(u24_16)) + -1.221268922091e-01*(V(u23_17) + V(u24_17))
+ + -1.944608241320e-01*(V(u23_18) + V(u24_18)) + -2.147991955280e-01*(V(u23_19) + V(u24_19)))
B_u32_2 u32_2 0 V = tanh_psi(2.114890813828e-01 + 1.673666238785e-01*(V(u23_0) + V(u24_0)) + -1.416311264038e-01*(V(u23_1) + V(u24_1))
+ + 2.127007544041e-01*(V(u23_2) + V(u24_2)) + -1.152877658606e-01*(V(u23_3) + V(u24_3)) + 9.290027618408e-02*(V(u23_4) + V(u24_4))
+ + -1.732315719128e-01*(V(u23_5) + V(u24_5)) + -7.225392758846e-02*(V(u23_6) + V(u24_6)) + 2.229158580303e-02*(V(u23_7) + V(u24_7))
+ + 8.696049451828e-03*(V(u23_8) + V(u24_8)) + -1.957250833511e-01*(V(u23_9) + V(u24_9)) + -2.387477457523e-02*(V(u23_10) + V(u24_10))
+ + -4.150708019733e-02*(V(u23_11) + V(u24_11)) + -2.033276855946e-01*(V(u23_12) + V(u24_12)) + 1.181437373161e-01*(V(u23_13)
+ + V(u24_13)) + 1.787683963776e-01*(V(u23_14) + V(u24_14)) + 1.052750349045e-01*(V(u23_15) + V(u24_15))
+ + 8.510792255402e-02*(V(u23_16) + V(u24_16)) + -8.157564699650e-02*(V(u23_17) + V(u24_17)) + -5.940197408199e-02*(V(u23_18)
+ + V(u24_18)) + 1.790322065353e-01*(V(u23_19) + V(u24_19)))
B_u32_3 u32_3 0 V = tanh_psi(7.760047912598e-02 + -2.121442109346e-01*(V(u23_0) + V(u24_0)) + 1.417499780655e-01*(V(u23_1) + V(u24_1))
+ + -1.688975244761e-01*(V(u23_2) + V(u24_2)) + -1.693129241467e-01*(V(u23_3) + V(u24_3)) + 1.521622836590e-01*(V(u23_4) + V(u24_4))
+ + -1.416471600533e-02*(V(u23_5) + V(u24_5)) + -1.168391704559e-01*(V(u23_6) + V(u24_6)) + -1.145977750421e-01*(V(u23_7) + V(u24_7))
+ + -1.938467770815e-01*(V(u23_8) + V(u24_8)) + -1.081197783351e-01*(V(u23_9) + V(u24_9)) + 1.430365145206e-01*(V(u23_10) + V(u24_10))
+ + -2.758646011353e-02*(V(u23_11) + V(u24_11)) + 1.033186912537e-02*(V(u23_12) + V(u24_12)) + -1.667422801256e-01*(V(u23_13)
+ + V(u24_13)) + 1.766636967659e-02*(V(u23_14) + V(u24_14)) + -1.971894949675e-01*(V(u23_15) + V(u24_15))
+ + 1.929947733879e-01*(V(u23_16) + V(u24_16)) + -1.720400154591e-02*(V(u23_17) + V(u24_17)) + 1.554751098156e-01*(V(u23_18)
+ + V(u24_18)) + -4.038918018341e-02*(V(u23_19) + V(u24_19)))
B_u32_4 u32_4 0 V = tanh_psi(3.173663020134e-01 + -1.783316731453e-01*(V(u23_0) + V(u24_0)) + -1.205225512385e-01*(V(u23_1) + V(u24_1))
+ + -1.368295848370e-01*(V(u23_2) + V(u24_2)) + 1.310324668884e-01*(V(u23_3) + V(u24_3)) + 1.065973937511e-02*(V(u23_4) + V(u24_4))
+ + 7.795971632004e-02*(V(u23_5) + V(u24_5)) + 1.457686126232e-01*(V(u23_6) + V(u24_6)) + 1.102370917797e-01*(V(u23_7) + V(u24_7))
+ + 5.112707614899e-03*(V(u23_8) + V(u24_8)) + -5.902814865112e-02*(V(u23_9) + V(u24_9)) + 2.122790217400e-01*(V(u23_10) + V(u24_10))
+ + -2.080718576908e-01*(V(u23_11) + V(u24_11)) + 1.162813901901e-01*(V(u23_12) + V(u24_12)) + 4.373431205750e-03*(V(u23_13)
+ + V(u24_13)) + -8.538654446602e-02*(V(u23_14) + V(u24_14)) + -2.831886708736e-02*(V(u23_15) + V(u24_15))
+ + 1.141825020313e-01*(V(u23_16) + V(u24_16)) + 7.949408888817e-02*(V(u23_17) + V(u24_17)) + -9.703859686852e-03*(V(u23_18)
+ + V(u24_18)) + -4.241800308228e-02*(V(u23_19) + V(u24_19)))
B_u32_5 u32_5 0 V = tanh_psi(1.712387204170e-01 + -1.871539652348e-02*(V(u23_0) + V(u24_0)) + 1.834868192673e-01*(V(u23_1) + V(u24_1))
+ + -2.049504369497e-01*(V(u23_2) + V(u24_2)) + 1.427587866783e-01*(V(u23_3) + V(u24_3)) + -2.132834494114e-02*(V(u23_4) + V(u24_4))
+ + -9.561800956726e-02*(V(u23_5) + V(u24_5)) + 2.144586741924e-01*(V(u23_6) + V(u24_6)) + 4.333209991455e-02*(V(u23_7) + V(u24_7))
+ + 1.173346340656e-01*(V(u23_8) + V(u24_8)) + 9.518310427666e-02*(V(u23_9) + V(u24_9)) + 1.481387019157e-01*(V(u23_10) + V(u24_10))
+ + -2.543911337852e-02*(V(u23_11) + V(u24_11)) + 6.930595636368e-02*(V(u23_12) + V(u24_12)) + 1.544605195522e-01*(V(u23_13)
+ + V(u24_13)) + -8.736599981785e-02*(V(u23_14) + V(u24_14)) + -4.072846472263e-02*(V(u23_15) + V(u24_15))
+ + 8.965235948563e-02*(V(u23_16) + V(u24_16)) + 8.628973364830e-02*(V(u23_17) + V(u24_17)) + 1.893289685249e-01*(V(u23_18)
+ + V(u24_18)) + -8.297756314278e-02*(V(u23_19) + V(u24_19)))
B_u32_6 u32_6 0 V = tanh_psi(-3.913363814354e-02 + -1.286404281855e-01*(V(u23_0) + V(u24_0)) + 1.118101775646e-01*(V(u23_1) + V(u24_1))
+ + -2.772240340710e-02*(V(u23_2) + V(u24_2)) + 3.766447305679e-03*(V(u23_3) + V(u24_3)) + -4.590477049351e-02*(V(u23_4) + V(u24_4))
+ + -7.390733063221e-02*(V(u23_5) + V(u24_5)) + -3.868146240711e-02*(V(u23_6) + V(u24_6)) + 5.403861403465e-02*(V(u23_7) + V(u24_7))
+ + 1.243321001530e-01*(V(u23_8) + V(u24_8)) + -2.349591255188e-02*(V(u23_9) + V(u24_9)) + -8.907006680965e-02*(V(u23_10) + V(u24_10))
+ + -1.105648502707e-01*(V(u23_11) + V(u24_11)) + -5.629138648510e-02*(V(u23_12) + V(u24_12)) + -1.420824825764e-01*(V(u23_13)
+ + V(u24_13)) + 6.944710016251e-02*(V(u23_14) + V(u24_14)) + -1.393491625786e-01*(V(u23_15) + V(u24_15))
+ + -7.176727056503e-02*(V(u23_16) + V(u24_16)) + 4.163280129433e-02*(V(u23_17) + V(u24_17)) + 1.304918229580e-01*(V(u23_18)
+ + V(u24_18)) + -1.462933123112e-01*(V(u23_19) + V(u24_19)))
B_u32_7 u32_7 0 V = tanh_psi(-3.302962481976e-01 + 1.531413197517e-01*(V(u23_0) + V(u24_0)) + 4.697009921074e-02*(V(u23_1) + V(u24_1))
+ + 8.314517140388e-02*(V(u23_2) + V(u24_2)) + 6.368109583855e-02*(V(u23_3) + V(u24_3)) + -1.248465478420e-02*(V(u23_4) + V(u24_4))
+ + -1.210482344031e-01*(V(u23_5) + V(u24_5)) + -8.373700082302e-02*(V(u23_6) + V(u24_6)) + 1.877845823765e-01*(V(u23_7) + V(u24_7))
+ + -2.812562882900e-02*(V(u23_8) + V(u24_8)) + -8.150026202202e-02*(V(u23_9) + V(u24_9)) + -1.647247374058e-02*(V(u23_10)
+ + V(u24_10)) + -8.729487657547e-02*(V(u23_11) + V(u24_11)) + -1.701740622520e-01*(V(u23_12) + V(u24_12))
+ + 4.201674461365e-02*(V(u23_13) + V(u24_13)) + -1.183368936181e-01*(V(u23_14) + V(u24_14)) + -1.012550592422e-01*(V(u23_15)
+ + V(u24_15)) + -1.535928547382e-01*(V(u23_16) + V(u24_16)) + 1.312710046768e-01*(V(u23_17) + V(u24_17))
+ + -7.475066184998e-02*(V(u23_18) + V(u24_18)) + -7.207331061363e-02*(V(u23_19) + V(u24_19)))
B_u32_8 u32_8 0 V = tanh_psi(1.790370941162e-01 + 2.384930849075e-04*(V(u23_0) + V(u24_0)) + -1.609933078289e-01*(V(u23_1) + V(u24_1))
+ + -8.743426203728e-02*(V(u23_2) + V(u24_2)) + -2.944640815258e-02*(V(u23_3) + V(u24_3)) + -1.944107413292e-01*(V(u23_4) + V(u24_4))
+ + -1.675792038441e-01*(V(u23_5) + V(u24_5)) + -3.022210299969e-02*(V(u23_6) + V(u24_6)) + 1.723698973656e-01*(V(u23_7) + V(u24_7))
+ + 1.015581786633e-01*(V(u23_8) + V(u24_8)) + 5.727520585060e-02*(V(u23_9) + V(u24_9)) + -6.700888276100e-03*(V(u23_10) + V(u24_10))
+ + -2.044115066528e-01*(V(u23_11) + V(u24_11)) + 1.579127907753e-01*(V(u23_12) + V(u24_12)) + 2.149165570736e-01*(V(u23_13)
+ + V(u24_13)) + 8.971634507179e-02*(V(u23_14) + V(u24_14)) + 1.126224398613e-01*(V(u23_15) + V(u24_15))
+ + -3.736537694931e-02*(V(u23_16) + V(u24_16)) + -1.748247593641e-01*(V(u23_17) + V(u24_17)) + -1.201171651483e-01*(V(u23_18)
+ + V(u24_18)) + 2.221004068851e-01*(V(u23_19) + V(u24_19)))
B_u32_9 u32_9 0 V = tanh_psi(-2.901732325554e-01 + 7.994458079338e-02*(V(u23_0) + V(u24_0)) + 1.125970780849e-01*(V(u23_1) + V(u24_1))
+ + -9.474912285805e-02*(V(u23_2) + V(u24_2)) + -1.131173223257e-01*(V(u23_3) + V(u24_3)) + 8.688080310822e-02*(V(u23_4) + V(u24_4))
+ + -1.801340430975e-01*(V(u23_5) + V(u24_5)) + 3.345751762390e-02*(V(u23_6) + V(u24_6)) + -1.838342845440e-02*(V(u23_7) + V(u24_7))
+ + 9.927454590797e-02*(V(u23_8) + V(u24_8)) + -1.252489089966e-01*(V(u23_9) + V(u24_9)) + 6.212249398232e-02*(V(u23_10) + V(u24_10))
+ + 4.049134254456e-02*(V(u23_11) + V(u24_11)) + -9.484082460403e-02*(V(u23_12) + V(u24_12)) + -1.879665702581e-01*(V(u23_13)
+ + V(u24_13)) + 7.639756798744e-02*(V(u23_14) + V(u24_14)) + -1.971459686756e-01*(V(u23_15) + V(u24_15))
+ + -9.454235434532e-02*(V(u23_16) + V(u24_16)) + -8.337506651878e-02*(V(u23_17) + V(u24_17)) + 1.742223203182e-01*(V(u23_18)
+ + V(u24_18)) + 2.597795426846e-02*(V(u23_19) + V(u24_19)))
B_u32_10 u32_10 0 V = tanh_psi(2.855592966080e-01 + -7.112193107605e-02*(V(u23_0) + V(u24_0)) + 1.412670314312e-02*(V(u23_1) + V(u24_1))
+ + 4.312169551849e-02*(V(u23_2) + V(u24_2)) + -3.987506031990e-03*(V(u23_3) + V(u24_3)) + 1.925032436848e-01*(V(u23_4) + V(u24_4))
+ + 1.595342755318e-01*(V(u23_5) + V(u24_5)) + -4.682341217995e-02*(V(u23_6) + V(u24_6)) + -7.670351862907e-02*(V(u23_7) + V(u24_7))
+ + -3.456015884876e-02*(V(u23_8) + V(u24_8)) + 5.525320768356e-02*(V(u23_9) + V(u24_9)) + -1.387401819229e-01*(V(u23_10) + V(u24_10))
+ + 1.947347223759e-01*(V(u23_11) + V(u24_11)) + 5.933240056038e-02*(V(u23_12) + V(u24_12)) + 1.615601778030e-01*(V(u23_13)
+ + V(u24_13)) + 1.002794802189e-01*(V(u23_14) + V(u24_14)) + -1.202769428492e-01*(V(u23_15) + V(u24_15))
+ + 8.291900157928e-04*(V(u23_16) + V(u24_16)) + -1.453912258148e-02*(V(u23_17) + V(u24_17)) + 1.802038848400e-01*(V(u23_18)
+ + V(u24_18)) + -1.447412073612e-01*(V(u23_19) + V(u24_19)))
B_u32_11 u32_11 0 V = tanh_psi(-1.133126020432e-02 + 1.357447803020e-01*(V(u23_0) + V(u24_0)) + -1.948305964470e-01*(V(u23_1) + V(u24_1))
+ + 5.361211299896e-02*(V(u23_2) + V(u24_2)) + -1.195701882243e-01*(V(u23_3) + V(u24_3)) + -2.431678771973e-02*(V(u23_4) + V(u24_4))
+ + -1.120856031775e-01*(V(u23_5) + V(u24_5)) + 5.906417965889e-03*(V(u23_6) + V(u24_6)) + 2.581439912319e-02*(V(u23_7) + V(u24_7))
+ + 9.321609139442e-02*(V(u23_8) + V(u24_8)) + -1.525077521801e-01*(V(u23_9) + V(u24_9)) + -1.121407747269e-02*(V(u23_10) + V(u24_10))
+ + 3.523662686348e-02*(V(u23_11) + V(u24_11)) + -4.172448813915e-02*(V(u23_12) + V(u24_12)) + 1.733103096485e-01*(V(u23_13)
+ + V(u24_13)) + 5.826562643051e-02*(V(u23_14) + V(u24_14)) + 2.217709124088e-01*(V(u23_15) + V(u24_15))
+ + -1.201465651393e-01*(V(u23_16) + V(u24_16)) + -5.016113817692e-02*(V(u23_17) + V(u24_17)) + -9.665286540985e-02*(V(u23_18)
+ + V(u24_18)) + 1.346867978573e-01*(V(u23_19) + V(u24_19)))
B_u32_12 u32_12 0 V = tanh_psi(-3.521715998650e-01 + 1.733688712120e-01*(V(u23_0) + V(u24_0)) + -7.884207367897e-02*(V(u23_1) + V(u24_1))
+ + -1.504434943199e-01*(V(u23_2) + V(u24_2)) + -8.206950128078e-02*(V(u23_3) + V(u24_3)) + 1.510509550571e-01*(V(u23_4) + V(u24_4))
+ + -1.439998298883e-01*(V(u23_5) + V(u24_5)) + -1.213082075119e-01*(V(u23_6) + V(u24_6)) + -1.998519748449e-01*(V(u23_7) + V(u24_7))
+ + 1.683471798897e-01*(V(u23_8) + V(u24_8)) + -1.158762499690e-01*(V(u23_9) + V(u24_9)) + -1.057954505086e-01*(V(u23_10) + V(u24_10))
+ + 1.220977604389e-01*(V(u23_11) + V(u24_11)) + -1.670566797256e-01*(V(u23_12) + V(u24_12)) + 1.242567896843e-01*(V(u23_13)
+ + V(u24_13)) + -1.174344494939e-01*(V(u23_14) + V(u24_14)) + -9.931457787752e-02*(V(u23_15) + V(u24_15))
+ + -3.638863563538e-05*(V(u23_16) + V(u24_16)) + 5.143147706985e-02*(V(u23_17) + V(u24_17)) + -1.699992716312e-01*(V(u23_18)
+ + V(u24_18)) + 9.619843959808e-02*(V(u23_19) + V(u24_19)))
B_u32_13 u32_13 0 V = tanh_psi(1.152889132500e-01 + -2.321565151215e-02*(V(u23_0) + V(u24_0)) + -1.857910901308e-01*(V(u23_1) + V(u24_1))
+ + 1.239010989666e-01*(V(u23_2) + V(u24_2)) + 1.184724569321e-01*(V(u23_3) + V(u24_3)) + -8.861760795116e-02*(V(u23_4) + V(u24_4))
+ + 1.141901314259e-01*(V(u23_5) + V(u24_5)) + 9.264451265335e-02*(V(u23_6) + V(u24_6)) + 1.798053383827e-01*(V(u23_7) + V(u24_7))
+ + 1.481645405293e-01*(V(u23_8) + V(u24_8)) + 3.749465942383e-02*(V(u23_9) + V(u24_9)) + 6.723478436470e-02*(V(u23_10) + V(u24_10))
+ + -1.723354607821e-01*(V(u23_11) + V(u24_11)) + -1.701672673225e-01*(V(u23_12) + V(u24_12)) + -1.267155408859e-01*(V(u23_13)
+ + V(u24_13)) + -1.762041449547e-02*(V(u23_14) + V(u24_14)) + -1.193560808897e-01*(V(u23_15) + V(u24_15))
+ + -1.760286390781e-01*(V(u23_16) + V(u24_16)) + -1.971642822027e-01*(V(u23_17) + V(u24_17)) + 1.317352652550e-01*(V(u23_18)
+ + V(u24_18)) + 1.364530324936e-01*(V(u23_19) + V(u24_19)))
B_u32_14 u32_14 0 V = tanh_psi(-2.415246963501e-01 + -1.479873806238e-01*(V(u23_0) + V(u24_0)) + 5.299851298332e-02*(V(u23_1) + V(u24_1))
+ + 5.294066667557e-02*(V(u23_2) + V(u24_2)) + 2.126453816891e-01*(V(u23_3) + V(u24_3)) + -2.166092991829e-01*(V(u23_4) + V(u24_4))
+ + -1.372461020947e-01*(V(u23_5) + V(u24_5)) + 4.980346560478e-02*(V(u23_6) + V(u24_6)) + 6.040748953819e-02*(V(u23_7) + V(u24_7))
+ + -8.354802429676e-02*(V(u23_8) + V(u24_8)) + -1.380520164967e-01*(V(u23_9) + V(u24_9)) + -6.867159903049e-02*(V(u23_10)
+ + V(u24_10)) + -5.551521480083e-02*(V(u23_11) + V(u24_11)) + -3.855139017105e-02*(V(u23_12) + V(u24_12))
+ + 6.145599484444e-02*(V(u23_13) + V(u24_13)) + -5.680991709232e-02*(V(u23_14) + V(u24_14)) + -8.434815704823e-02*(V(u23_15)
+ + V(u24_15)) + -1.199336126447e-01*(V(u23_16) + V(u24_16)) + 7.883039116859e-02*(V(u23_17) + V(u24_17))
+ + -7.586456835270e-02*(V(u23_18) + V(u24_18)) + -6.863473355770e-02*(V(u23_19) + V(u24_19)))
B_u32_15 u32_15 0 V = tanh_psi(1.432535648346e-01 + -1.773540675640e-01*(V(u23_0) + V(u24_0)) + -1.086149960756e-01*(V(u23_1) + V(u24_1))
+ + -5.619721114635e-02*(V(u23_2) + V(u24_2)) + -8.678416907787e-02*(V(u23_3) + V(u24_3)) + -2.168527692556e-01*(V(u23_4) + V(u24_4))
+ + -4.911760985851e-02*(V(u23_5) + V(u24_5)) + 1.907641589642e-01*(V(u23_6) + V(u24_6)) + -1.908497661352e-01*(V(u23_7) + V(u24_7))
+ + -1.274053156376e-01*(V(u23_8) + V(u24_8)) + 5.828055739403e-02*(V(u23_9) + V(u24_9)) + 2.167389094830e-01*(V(u23_10) + V(u24_10))
+ + 2.068177759647e-01*(V(u23_11) + V(u24_11)) + -3.971262276173e-02*(V(u23_12) + V(u24_12)) + -1.836395263672e-01*(V(u23_13)
+ + V(u24_13)) + 1.841551065445e-01*(V(u23_14) + V(u24_14)) + 2.078063189983e-01*(V(u23_15) + V(u24_15))
+ + 1.238479018211e-01*(V(u23_16) + V(u24_16)) + 1.209149956703e-01*(V(u23_17) + V(u24_17)) + 1.189693808556e-01*(V(u23_18)
+ + V(u24_18)) + -1.121744737029e-01*(V(u23_19) + V(u24_19)))
B_u32_16 u32_16 0 V = tanh_psi(-4.338133335114e-02 + -1.844362765551e-01*(V(u23_0) + V(u24_0)) + 1.900017857552e-01*(V(u23_1) + V(u24_1))
+ + 2.119104862213e-01*(V(u23_2) + V(u24_2)) + 1.628711223602e-01*(V(u23_3) + V(u24_3)) + -2.159997522831e-01*(V(u23_4) + V(u24_4))
+ + 1.250273883343e-01*(V(u23_5) + V(u24_5)) + -1.784750819206e-01*(V(u23_6) + V(u24_6)) + -4.456785321236e-02*(V(u23_7) + V(u24_7))
+ + 2.219927608967e-01*(V(u23_8) + V(u24_8)) + -9.556381404400e-02*(V(u23_9) + V(u24_9)) + 1.063317358494e-01*(V(u23_10) + V(u24_10))
+ + 1.297687888145e-01*(V(u23_11) + V(u24_11)) + -6.874610483646e-02*(V(u23_12) + V(u24_12)) + 2.165578603745e-01*(V(u23_13)
+ + V(u24_13)) + 2.087486088276e-01*(V(u23_14) + V(u24_14)) + 1.043610274792e-01*(V(u23_15) + V(u24_15))
+ + -5.802474915981e-02*(V(u23_16) + V(u24_16)) + -1.534143835306e-01*(V(u23_17) + V(u24_17)) + 1.827417910099e-01*(V(u23_18)
+ + V(u24_18)) + -2.124366164207e-02*(V(u23_19) + V(u24_19)))
B_u32_17 u32_17 0 V = tanh_psi(-1.626423597336e-01 + -1.423172652721e-02*(V(u23_0) + V(u24_0)) + 1.306897699833e-01*(V(u23_1) + V(u24_1))
+ + -1.327999085188e-01*(V(u23_2) + V(u24_2)) + 2.224712371826e-01*(V(u23_3) + V(u24_3)) + -5.315743386745e-02*(V(u23_4) + V(u24_4))
+ + 1.119352877140e-02*(V(u23_5) + V(u24_5)) + 2.102293968201e-01*(V(u23_6) + V(u24_6)) + 1.594474017620e-01*(V(u23_7) + V(u24_7))
+ + 8.160710334778e-02*(V(u23_8) + V(u24_8)) + -2.215330302715e-01*(V(u23_9) + V(u24_9)) + 1.335639357567e-01*(V(u23_10) + V(u24_10))
+ + 1.401656866074e-01*(V(u23_11) + V(u24_11)) + -3.000080585480e-03*(V(u23_12) + V(u24_12)) + 1.916750371456e-01*(V(u23_13)
+ + V(u24_13)) + 1.075125038624e-01*(V(u23_14) + V(u24_14)) + 1.173050403595e-01*(V(u23_15) + V(u24_15))
+ + 1.030759513378e-01*(V(u23_16) + V(u24_16)) + -1.027870550752e-01*(V(u23_17) + V(u24_17)) + -2.781556546688e-02*(V(u23_18)
+ + V(u24_18)) + -2.206156700850e-01*(V(u23_19) + V(u24_19)))
B_u32_18 u32_18 0 V = tanh_psi(-2.598097026348e-01 + -2.020823657513e-01*(V(u23_0) + V(u24_0)) + -1.912469118834e-01*(V(u23_1) + V(u24_1))
+ + 1.209463179111e-01*(V(u23_2) + V(u24_2)) + 1.091353297234e-01*(V(u23_3) + V(u24_3)) + 1.627348065376e-01*(V(u23_4) + V(u24_4))
+ + 2.156421244144e-01*(V(u23_5) + V(u24_5)) + -2.184545695782e-01*(V(u23_6) + V(u24_6)) + 2.357637882233e-02*(V(u23_7) + V(u24_7))
+ + 2.155182659626e-01*(V(u23_8) + V(u24_8)) + -3.467938303947e-02*(V(u23_9) + V(u24_9)) + -1.414653658867e-02*(V(u23_10) + V(u24_10))
+ + -6.224191188812e-02*(V(u23_11) + V(u24_11)) + -7.254709303379e-02*(V(u23_12) + V(u24_12)) + 1.407925486565e-01*(V(u23_13)
+ + V(u24_13)) + 1.526156663895e-01*(V(u23_14) + V(u24_14)) + -1.460507512093e-01*(V(u23_15) + V(u24_15))
+ + -1.763346642256e-01*(V(u23_16) + V(u24_16)) + 2.163420617580e-01*(V(u23_17) + V(u24_17)) + 1.481215655804e-01*(V(u23_18)
+ + V(u24_18)) + 1.975628733635e-02*(V(u23_19) + V(u24_19)))
B_u32_19 u32_19 0 V = tanh_psi(2.660924196243e-01 + -2.043821066618e-01*(V(u23_0) + V(u24_0)) + 1.583797931671e-01*(V(u23_1) + V(u24_1))
+ + -1.807579547167e-01*(V(u23_2) + V(u24_2)) + -1.904599964619e-01*(V(u23_3) + V(u24_3)) + 1.426028609276e-01*(V(u23_4) + V(u24_4))
+ + 2.038039267063e-01*(V(u23_5) + V(u24_5)) + 7.856833934784e-02*(V(u23_6) + V(u24_6)) + 6.092542409897e-02*(V(u23_7) + V(u24_7))
+ + -1.601629108191e-01*(V(u23_8) + V(u24_8)) + 1.971647441387e-01*(V(u23_9) + V(u24_9)) + -1.547144353390e-01*(V(u23_10) + V(u24_10))
+ + 1.914219558239e-01*(V(u23_11) + V(u24_11)) + -2.790844440460e-02*(V(u23_12) + V(u24_12)) + 2.967157959938e-02*(V(u23_13)
+ + V(u24_13)) + -6.683005392551e-02*(V(u23_14) + V(u24_14)) + -1.089076772332e-01*(V(u23_15) + V(u24_15))
+ + -1.494662314653e-01*(V(u23_16) + V(u24_16)) + 7.819998264313e-02*(V(u23_17) + V(u24_17)) + -2.282233536243e-02*(V(u23_18)
+ + V(u24_18)) + 1.433448195457e-01*(V(u23_19) + V(u24_19)))
B_u32_20 u32_20 0 V = tanh_psi(-3.214898407459e-01 + 1.604641377926e-01*(V(u23_0) + V(u24_0)) + -1.651054471731e-01*(V(u23_1) + V(u24_1))
+ + -4.967102408409e-02*(V(u23_2) + V(u24_2)) + -1.665388196707e-01*(V(u23_3) + V(u24_3)) + 5.796256661415e-02*(V(u23_4) + V(u24_4))
+ + -1.019986495376e-01*(V(u23_5) + V(u24_5)) + 1.522459089756e-01*(V(u23_6) + V(u24_6)) + 6.798979640007e-02*(V(u23_7) + V(u24_7))
+ + -1.407386958599e-01*(V(u23_8) + V(u24_8)) + -1.453046202660e-01*(V(u23_9) + V(u24_9)) + 1.237377524376e-03*(V(u23_10) + V(u24_10))
+ + 1.613025367260e-01*(V(u23_11) + V(u24_11)) + -9.402424097061e-03*(V(u23_12) + V(u24_12)) + -2.018473595381e-01*(V(u23_13)
+ + V(u24_13)) + -1.339356601238e-01*(V(u23_14) + V(u24_14)) + -8.522252738476e-02*(V(u23_15) + V(u24_15))
+ + -2.081535607576e-01*(V(u23_16) + V(u24_16)) + -1.141830310225e-01*(V(u23_17) + V(u24_17)) + -2.015406042337e-01*(V(u23_18)
+ + V(u24_18)) + -1.369178295135e-01*(V(u23_19) + V(u24_19)))
B_u32_21 u32_21 0 V = tanh_psi(-4.421823620796e-01 + 1.051650941372e-02*(V(u23_0) + V(u24_0)) + 3.242895007133e-03*(V(u23_1) + V(u24_1))
+ + 4.978761076927e-02*(V(u23_2) + V(u24_2)) + 9.213060140610e-02*(V(u23_3) + V(u24_3)) + 1.033160090446e-01*(V(u23_4) + V(u24_4))
+ + 2.023664712906e-01*(V(u23_5) + V(u24_5)) + 9.179183840752e-02*(V(u23_6) + V(u24_6)) + 1.656068861485e-02*(V(u23_7) + V(u24_7))
+ + -1.325068175793e-01*(V(u23_8) + V(u24_8)) + 1.176698803902e-01*(V(u23_9) + V(u24_9)) + -1.076386347413e-01*(V(u23_10) + V(u24_10))
+ + 7.383203506470e-02*(V(u23_11) + V(u24_11)) + -7.898376882076e-02*(V(u23_12) + V(u24_12)) + -1.119541078806e-01*(V(u23_13)
+ + V(u24_13)) + 1.908402740955e-01*(V(u23_14) + V(u24_14)) + -2.179072648287e-01*(V(u23_15) + V(u24_15))
+ + 1.322558224201e-01*(V(u23_16) + V(u24_16)) + 5.072921514511e-02*(V(u23_17) + V(u24_17)) + 1.921981275082e-01*(V(u23_18)
+ + V(u24_18)) + -5.215439200401e-02*(V(u23_19) + V(u24_19)))
B_u32_22 u32_22 0 V = tanh_psi(-4.239812791348e-01 + -2.206100225449e-01*(V(u23_0) + V(u24_0)) + 8.456316590309e-02*(V(u23_1) + V(u24_1))
+ + 1.504628360271e-02*(V(u23_2) + V(u24_2)) + 5.737441778183e-02*(V(u23_3) + V(u24_3)) + -1.585682183504e-01*(V(u23_4) + V(u24_4))
+ + 4.794076085091e-02*(V(u23_5) + V(u24_5)) + -5.418919026852e-02*(V(u23_6) + V(u24_6)) + -1.988849192858e-01*(V(u23_7) + V(u24_7))
+ + -1.245507523417e-01*(V(u23_8) + V(u24_8)) + 1.112564504147e-01*(V(u23_9) + V(u24_9)) + 1.841324269772e-01*(V(u23_10) + V(u24_10))
+ + 1.252453923225e-01*(V(u23_11) + V(u24_11)) + -1.711940765381e-01*(V(u23_12) + V(u24_12)) + 5.306944251060e-02*(V(u23_13)
+ + V(u24_13)) + 5.557367205620e-02*(V(u23_14) + V(u24_14)) + 2.226187288761e-01*(V(u23_15) + V(u24_15))
+ + -6.926774978638e-03*(V(u23_16) + V(u24_16)) + 1.675815284252e-01*(V(u23_17) + V(u24_17)) + -5.505184829235e-02*(V(u23_18)
+ + V(u24_18)) + -1.105124205351e-01*(V(u23_19) + V(u24_19)))
B_u32_23 u32_23 0 V = tanh_psi(-2.985839545727e-01 + -1.570796370506e-01*(V(u23_0) + V(u24_0)) + -6.177966296673e-02*(V(u23_1) + V(u24_1))
+ + 2.078866362572e-01*(V(u23_2) + V(u24_2)) + 5.788356065750e-02*(V(u23_3) + V(u24_3)) + 1.233199536800e-01*(V(u23_4) + V(u24_4))
+ + 1.099173128605e-01*(V(u23_5) + V(u24_5)) + 1.974871754646e-02*(V(u23_6) + V(u24_6)) + 8.757692575455e-02*(V(u23_7) + V(u24_7))
+ + -1.072780042887e-01*(V(u23_8) + V(u24_8)) + -1.538584828377e-01*(V(u23_9) + V(u24_9)) + 1.702217161655e-01*(V(u23_10) + V(u24_10))
+ + -1.126601994038e-01*(V(u23_11) + V(u24_11)) + -6.260165572166e-02*(V(u23_12) + V(u24_12)) + 1.878895461559e-01*(V(u23_13)
+ + V(u24_13)) + -9.866657108068e-02*(V(u23_14) + V(u24_14)) + -2.080154567957e-01*(V(u23_15) + V(u24_15))
+ + 1.047514677048e-01*(V(u23_16) + V(u24_16)) + -2.130653560162e-01*(V(u23_17) + V(u24_17)) + -1.060148030519e-01*(V(u23_18)
+ + V(u24_18)) + -1.304394900799e-01*(V(u23_19) + V(u24_19)))
B_u32_24 u32_24 0 V = tanh_psi(-3.199982047081e-01 + -1.862553060055e-01*(V(u23_0) + V(u24_0)) + 4.422485828400e-02*(V(u23_1) + V(u24_1))
+ + -2.232264727354e-01*(V(u23_2) + V(u24_2)) + -1.032869666815e-01*(V(u23_3) + V(u24_3)) + 1.262583136559e-01*(V(u23_4) + V(u24_4))
+ + -3.445845842361e-02*(V(u23_5) + V(u24_5)) + -5.855183303356e-02*(V(u23_6) + V(u24_6)) + -1.950900107622e-01*(V(u23_7) + V(u24_7))
+ + 2.149181365967e-01*(V(u23_8) + V(u24_8)) + -1.367225497961e-01*(V(u23_9) + V(u24_9)) + 2.057889401913e-01*(V(u23_10) + V(u24_10))
+ + -5.543388426304e-02*(V(u23_11) + V(u24_11)) + 8.573451638222e-02*(V(u23_12) + V(u24_12)) + -5.054591596127e-02*(V(u23_13)
+ + V(u24_13)) + 1.445088386536e-01*(V(u23_14) + V(u24_14)) + 3.823995590210e-03*(V(u23_15) + V(u24_15))
+ + -1.345014870167e-01*(V(u23_16) + V(u24_16)) + -1.316874176264e-01*(V(u23_17) + V(u24_17)) + 7.119065523148e-02*(V(u23_18)
+ + V(u24_18)) + -7.532036304474e-02*(V(u23_19) + V(u24_19)))
B_u32_25 u32_25 0 V = tanh_psi(2.934380173683e-01 + 1.431837677956e-01*(V(u23_0) + V(u24_0)) + 1.862487196922e-01*(V(u23_1) + V(u24_1))
+ + 1.851477921009e-01*(V(u23_2) + V(u24_2)) + 8.680829405785e-02*(V(u23_3) + V(u24_3)) + 6.356501579285e-02*(V(u23_4) + V(u24_4))
+ + 1.759128570557e-01*(V(u23_5) + V(u24_5)) + -1.884937286377e-02*(V(u23_6) + V(u24_6)) + -1.064942106605e-01*(V(u23_7) + V(u24_7))
+ + -2.133840024471e-01*(V(u23_8) + V(u24_8)) + 1.061036884785e-01*(V(u23_9) + V(u24_9)) + 1.447155475616e-01*(V(u23_10) + V(u24_10))
+ + 7.768628001213e-02*(V(u23_11) + V(u24_11)) + -4.484950006008e-02*(V(u23_12) + V(u24_12)) + -8.129112422466e-02*(V(u23_13)
+ + V(u24_13)) + -2.096398472786e-01*(V(u23_14) + V(u24_14)) + -1.791086494923e-01*(V(u23_15) + V(u24_15))
+ + -1.210442632437e-01*(V(u23_16) + V(u24_16)) + -2.031293362379e-01*(V(u23_17) + V(u24_17)) + 9.447771310806e-02*(V(u23_18)
+ + V(u24_18)) + -1.516643166542e-01*(V(u23_19) + V(u24_19)))
B_u32_26 u32_26 0 V = tanh_psi(-9.157085418701e-02 + -1.189523935318e-02*(V(u23_0) + V(u24_0)) + -1.046681478620e-01*(V(u23_1) + V(u24_1))
+ + -4.573406279087e-02*(V(u23_2) + V(u24_2)) + 4.577720165253e-02*(V(u23_3) + V(u24_3)) + -3.008238971233e-02*(V(u23_4) + V(u24_4))
+ + -4.572777450085e-02*(V(u23_5) + V(u24_5)) + -1.810698807240e-01*(V(u23_6) + V(u24_6)) + 5.750244855881e-02*(V(u23_7) + V(u24_7))
+ + 2.091141939163e-01*(V(u23_8) + V(u24_8)) + -1.483143866062e-01*(V(u23_9) + V(u24_9)) + 3.725728392601e-02*(V(u23_10) + V(u24_10))
+ + -1.568057239056e-01*(V(u23_11) + V(u24_11)) + -2.217176854610e-01*(V(u23_12) + V(u24_12)) + -3.930652141571e-02*(V(u23_13)
+ + V(u24_13)) + -1.654887795448e-01*(V(u23_14) + V(u24_14)) + -1.253442466259e-02*(V(u23_15) + V(u24_15))
+ + -2.112434208393e-01*(V(u23_16) + V(u24_16)) + -3.055720031261e-02*(V(u23_17) + V(u24_17)) + 9.331557154655e-02*(V(u23_18)
+ + V(u24_18)) + 3.279379010201e-02*(V(u23_19) + V(u24_19)))
B_u32_27 u32_27 0 V = tanh_psi(2.278879284859e-01 + -1.522485911846e-01*(V(u23_0) + V(u24_0)) + -1.341211497784e-01*(V(u23_1) + V(u24_1))
+ + -1.661857068539e-01*(V(u23_2) + V(u24_2)) + -9.302373230457e-02*(V(u23_3) + V(u24_3)) + 1.669228374958e-01*(V(u23_4) + V(u24_4))
+ + -7.304905354977e-02*(V(u23_5) + V(u24_5)) + -8.627611398697e-02*(V(u23_6) + V(u24_6)) + -1.578655391932e-01*(V(u23_7) + V(u24_7))
+ + 1.622292399406e-01*(V(u23_8) + V(u24_8)) + 1.071792244911e-01*(V(u23_9) + V(u24_9)) + 9.333443641663e-02*(V(u23_10) + V(u24_10))
+ + 2.160333395004e-01*(V(u23_11) + V(u24_11)) + -1.879915446043e-01*(V(u23_12) + V(u24_12)) + -5.165526270866e-02*(V(u23_13)
+ + V(u24_13)) + 2.084893584251e-01*(V(u23_14) + V(u24_14)) + -7.990959286690e-02*(V(u23_15) + V(u24_15))
+ + 5.936628580093e-02*(V(u23_16) + V(u24_16)) + -4.756610095501e-02*(V(u23_17) + V(u24_17)) + -4.466570913792e-02*(V(u23_18)
+ + V(u24_18)) + 1.501283943653e-01*(V(u23_19) + V(u24_19)))
B_u32_28 u32_28 0 V = tanh_psi(-6.358012557030e-02 + -2.122449874878e-01*(V(u23_0) + V(u24_0)) + -1.353091746569e-01*(V(u23_1) + V(u24_1))
+ + -1.033015474677e-01*(V(u23_2) + V(u24_2)) + 2.694860100746e-02*(V(u23_3) + V(u24_3)) + -1.590049564838e-01*(V(u23_4) + V(u24_4))
+ + 1.420590281487e-01*(V(u23_5) + V(u24_5)) + 2.153514325619e-02*(V(u23_6) + V(u24_6)) + 6.975471973419e-02*(V(u23_7) + V(u24_7))
+ + -1.955806463957e-01*(V(u23_8) + V(u24_8)) + 7.233941555023e-02*(V(u23_9) + V(u24_9)) + 1.943807303905e-01*(V(u23_10) + V(u24_10))
+ + -1.061895340681e-01*(V(u23_11) + V(u24_11)) + 1.917980313301e-01*(V(u23_12) + V(u24_12)) + -1.914220899343e-01*(V(u23_13)
+ + V(u24_13)) + -2.025910913944e-01*(V(u23_14) + V(u24_14)) + -1.231198087335e-01*(V(u23_15) + V(u24_15))
+ + -1.656920909882e-01*(V(u23_16) + V(u24_16)) + -1.455669105053e-02*(V(u23_17) + V(u24_17)) + -1.693422496319e-01*(V(u23_18)
+ + V(u24_18)) + -1.968954503536e-01*(V(u23_19) + V(u24_19)))
B_u32_29 u32_29 0 V = tanh_psi(3.906453251839e-01 + -9.149122238159e-02*(V(u23_0) + V(u24_0)) + 1.705335676670e-01*(V(u23_1) + V(u24_1))
+ + 1.600608229637e-02*(V(u23_2) + V(u24_2)) + -1.425226926804e-01*(V(u23_3) + V(u24_3)) + -4.444727301598e-02*(V(u23_4) + V(u24_4))
+ + -1.055138036609e-01*(V(u23_5) + V(u24_5)) + -8.730199933052e-02*(V(u23_6) + V(u24_6)) + -9.471130371094e-02*(V(u23_7) + V(u24_7))
+ + -1.171212419868e-01*(V(u23_8) + V(u24_8)) + -1.835702955723e-01*(V(u23_9) + V(u24_9)) + 5.953520536423e-02*(V(u23_10) + V(u24_10))
+ + -2.118215560913e-01*(V(u23_11) + V(u24_11)) + 2.523796260357e-02*(V(u23_12) + V(u24_12)) + 5.455499887466e-02*(V(u23_13)
+ + V(u24_13)) + -1.573662161827e-01*(V(u23_14) + V(u24_14)) + -1.056749448180e-01*(V(u23_15) + V(u24_15))
+ + 1.155340671539e-02*(V(u23_16) + V(u24_16)) + 1.258700191975e-01*(V(u23_17) + V(u24_17)) + 1.117213964462e-01*(V(u23_18)
+ + V(u24_18)) + -1.183973178267e-01*(V(u23_19) + V(u24_19)))
B_u32_30 u32_30 0 V = tanh_psi(-4.838779568672e-02 + -1.211600303650e-01*(V(u23_0) + V(u24_0)) + 1.666389405727e-01*(V(u23_1) + V(u24_1))
+ + -3.276795148849e-03*(V(u23_2) + V(u24_2)) + -8.047835528851e-02*(V(u23_3) + V(u24_3)) + 2.004212737083e-01*(V(u23_4) + V(u24_4))
+ + -1.789529770613e-01*(V(u23_5) + V(u24_5)) + -2.045704424381e-02*(V(u23_6) + V(u24_6)) + 7.913088798523e-02*(V(u23_7) + V(u24_7))
+ + -1.036944538355e-01*(V(u23_8) + V(u24_8)) + 2.630892395973e-02*(V(u23_9) + V(u24_9)) + -2.118208408356e-01*(V(u23_10) + V(u24_10))
+ + -1.232836619020e-01*(V(u23_11) + V(u24_11)) + -1.425628811121e-01*(V(u23_12) + V(u24_12)) + 1.940868198872e-01*(V(u23_13)
+ + V(u24_13)) + 2.226270139217e-01*(V(u23_14) + V(u24_14)) + 1.283576488495e-01*(V(u23_15) + V(u24_15))
+ + 1.818298995495e-01*(V(u23_16) + V(u24_16)) + 8.874937891960e-02*(V(u23_17) + V(u24_17)) + -6.296470761299e-03*(V(u23_18)
+ + V(u24_18)) + -3.225998580456e-02*(V(u23_19) + V(u24_19)))
B_u32_31 u32_31 0 V = tanh_psi(7.532590627670e-02 + 1.718633472919e-01*(V(u23_0) + V(u24_0)) + -4.762105643749e-02*(V(u23_1) + V(u24_1))
+ + -1.257322728634e-01*(V(u23_2) + V(u24_2)) + 1.397567391396e-01*(V(u23_3) + V(u24_3)) + 5.273637175560e-02*(V(u23_4) + V(u24_4))
+ + 1.483164131641e-01*(V(u23_5) + V(u24_5)) + -1.199399605393e-01*(V(u23_6) + V(u24_6)) + 1.137101948261e-01*(V(u23_7) + V(u24_7))
+ + -1.061810329556e-01*(V(u23_8) + V(u24_8)) + 1.761509180069e-01*(V(u23_9) + V(u24_9)) + 2.306294441223e-02*(V(u23_10) + V(u24_10))
+ + -7.840481400490e-02*(V(u23_11) + V(u24_11)) + -9.979982674122e-02*(V(u23_12) + V(u24_12)) + -1.014747843146e-01*(V(u23_13)
+ + V(u24_13)) + -1.868531703949e-01*(V(u23_14) + V(u24_14)) + 4.937201738358e-03*(V(u23_15) + V(u24_15))
+ + 5.807110667229e-02*(V(u23_16) + V(u24_16)) + -1.423737853765e-01*(V(u23_17) + V(u24_17)) + 8.230715990067e-03*(V(u23_18)
+ + V(u24_18)) + 1.142345368862e-01*(V(u23_19) + V(u24_19)))
B_u32_32 u32_32 0 V = tanh_psi(6.743037700653e-02 + 1.348994076252e-01*(V(u23_0) + V(u24_0)) + -1.863270848989e-01*(V(u23_1) + V(u24_1))
+ + -3.842404484749e-02*(V(u23_2) + V(u24_2)) + 7.793602347374e-02*(V(u23_3) + V(u24_3)) + 1.917437314987e-01*(V(u23_4) + V(u24_4))
+ + -7.213155925274e-02*(V(u23_5) + V(u24_5)) + 1.605929434299e-01*(V(u23_6) + V(u24_6)) + 5.562993884087e-02*(V(u23_7) + V(u24_7))
+ + 1.418458819389e-01*(V(u23_8) + V(u24_8)) + 1.065450608730e-01*(V(u23_9) + V(u24_9)) + -8.796642720699e-02*(V(u23_10) + V(u24_10))
+ + 1.181851625443e-01*(V(u23_11) + V(u24_11)) + 1.199119985104e-01*(V(u23_12) + V(u24_12)) + 2.172632515430e-02*(V(u23_13)
+ + V(u24_13)) + 2.110709547997e-01*(V(u23_14) + V(u24_14)) + -1.344622373581e-01*(V(u23_15) + V(u24_15))
+ + 1.029575169086e-01*(V(u23_16) + V(u24_16)) + -1.693892478943e-01*(V(u23_17) + V(u24_17)) + 2.079021036625e-01*(V(u23_18)
+ + V(u24_18)) + -4.619246721268e-02*(V(u23_19) + V(u24_19)))
B_u32_33 u32_33 0 V = tanh_psi(-2.627612650394e-01 + -1.924925446510e-01*(V(u23_0) + V(u24_0)) + 2.025640010834e-02*(V(u23_1) + V(u24_1))
+ + -1.264923810959e-01*(V(u23_2) + V(u24_2)) + -1.360898166895e-01*(V(u23_3) + V(u24_3)) + -8.268462121487e-02*(V(u23_4) + V(u24_4))
+ + -4.781568050385e-02*(V(u23_5) + V(u24_5)) + -1.410123556852e-01*(V(u23_6) + V(u24_6)) + -1.719504147768e-01*(V(u23_7) + V(u24_7))
+ + 1.028715670109e-01*(V(u23_8) + V(u24_8)) + 1.443094313145e-01*(V(u23_9) + V(u24_9)) + 8.423456549644e-02*(V(u23_10) + V(u24_10))
+ + 1.135935783386e-01*(V(u23_11) + V(u24_11)) + -1.567694693804e-01*(V(u23_12) + V(u24_12)) + 5.035474896431e-03*(V(u23_13)
+ + V(u24_13)) + 2.634325623512e-02*(V(u23_14) + V(u24_14)) + -1.910185515881e-01*(V(u23_15) + V(u24_15))
+ + 6.578016281128e-02*(V(u23_16) + V(u24_16)) + 6.787255406380e-03*(V(u23_17) + V(u24_17)) + -5.784361064434e-02*(V(u23_18)
+ + V(u24_18)) + 9.846994280815e-02*(V(u23_19) + V(u24_19)))
B_u32_34 u32_34 0 V = tanh_psi(-2.755779027939e-01 + 1.849233210087e-01*(V(u23_0) + V(u24_0)) + 7.098788022995e-02*(V(u23_1) + V(u24_1))
+ + -1.717496663332e-01*(V(u23_2) + V(u24_2)) + 1.908898353577e-02*(V(u23_3) + V(u24_3)) + -7.912401854992e-02*(V(u23_4) + V(u24_4))
+ + 2.116540074348e-01*(V(u23_5) + V(u24_5)) + -2.144017815590e-02*(V(u23_6) + V(u24_6)) + 1.483735144138e-01*(V(u23_7) + V(u24_7))
+ + 4.250967502594e-02*(V(u23_8) + V(u24_8)) + 2.189510166645e-01*(V(u23_9) + V(u24_9)) + -2.305662631989e-02*(V(u23_10) + V(u24_10))
+ + 4.206931591034e-02*(V(u23_11) + V(u24_11)) + -1.243998110294e-02*(V(u23_12) + V(u24_12)) + 1.084871888161e-01*(V(u23_13)
+ + V(u24_13)) + -4.942898452282e-02*(V(u23_14) + V(u24_14)) + -1.880155056715e-01*(V(u23_15) + V(u24_15))
+ + 5.870571732521e-02*(V(u23_16) + V(u24_16)) + -2.026848196983e-01*(V(u23_17) + V(u24_17)) + -4.734413325787e-02*(V(u23_18)
+ + V(u24_18)) + 9.014013409615e-02*(V(u23_19) + V(u24_19)))
B_u32_35 u32_35 0 V = tanh_psi(2.275888323784e-01 + 2.088822722435e-01*(V(u23_0) + V(u24_0)) + 2.012824714184e-01*(V(u23_1) + V(u24_1))
+ + 1.302275955677e-01*(V(u23_2) + V(u24_2)) + -5.293981730938e-02*(V(u23_3) + V(u24_3)) + 1.928474605083e-01*(V(u23_4) + V(u24_4))
+ + 4.249259829521e-03*(V(u23_5) + V(u24_5)) + 1.981941163540e-01*(V(u23_6) + V(u24_6)) + 2.010024487972e-01*(V(u23_7) + V(u24_7))
+ + 1.310379207134e-01*(V(u23_8) + V(u24_8)) + 1.461072266102e-01*(V(u23_9) + V(u24_9)) + 1.334953904152e-01*(V(u23_10) + V(u24_10))
+ + -2.920219302177e-02*(V(u23_11) + V(u24_11)) + -1.097046136856e-01*(V(u23_12) + V(u24_12)) + -1.524068713188e-01*(V(u23_13)
+ + V(u24_13)) + 2.069935798645e-01*(V(u23_14) + V(u24_14)) + 4.110002517700e-02*(V(u23_15) + V(u24_15))
+ + -3.433480858803e-02*(V(u23_16) + V(u24_16)) + 7.806688547134e-02*(V(u23_17) + V(u24_17)) + 1.713167428970e-01*(V(u23_18)
+ + V(u24_18)) + -9.988973289728e-02*(V(u23_19) + V(u24_19)))
B_u32_36 u32_36 0 V = tanh_psi(-2.301891297102e-01 + 2.180243432522e-01*(V(u23_0) + V(u24_0)) + 9.238103032112e-02*(V(u23_1) + V(u24_1))
+ + -2.128224968910e-01*(V(u23_2) + V(u24_2)) + 2.861350774765e-02*(V(u23_3) + V(u24_3)) + -6.966227293015e-02*(V(u23_4) + V(u24_4))
+ + 1.830382049084e-01*(V(u23_5) + V(u24_5)) + 1.798828244209e-01*(V(u23_6) + V(u24_6)) + -1.422844529152e-01*(V(u23_7) + V(u24_7))
+ + 1.707144379616e-01*(V(u23_8) + V(u24_8)) + -4.939630627632e-02*(V(u23_9) + V(u24_9)) + 1.659149825573e-01*(V(u23_10) + V(u24_10))
+ + -4.155918955803e-02*(V(u23_11) + V(u24_11)) + -7.802200317383e-02*(V(u23_12) + V(u24_12)) + 1.695597767830e-01*(V(u23_13)
+ + V(u24_13)) + -6.372012197971e-02*(V(u23_14) + V(u24_14)) + 1.208730041981e-01*(V(u23_15) + V(u24_15))
+ + 1.185298264027e-01*(V(u23_16) + V(u24_16)) + 9.795612096786e-02*(V(u23_17) + V(u24_17)) + 1.430476009846e-01*(V(u23_18)
+ + V(u24_18)) + 2.172589302063e-05*(V(u23_19) + V(u24_19)))
B_u32_37 u32_37 0 V = tanh_psi(-2.902398705482e-01 + -9.104415774345e-02*(V(u23_0) + V(u24_0)) + 9.930178523064e-02*(V(u23_1) + V(u24_1))
+ + -1.405076980591e-01*(V(u23_2) + V(u24_2)) + -1.053378731012e-01*(V(u23_3) + V(u24_3)) + 5.724072456360e-02*(V(u23_4) + V(u24_4))
+ + -5.107024312019e-02*(V(u23_5) + V(u24_5)) + -1.459648311138e-01*(V(u23_6) + V(u24_6)) + -1.988439261913e-01*(V(u23_7) + V(u24_7))
+ + 8.278346061707e-02*(V(u23_8) + V(u24_8)) + -1.662615686655e-01*(V(u23_9) + V(u24_9)) + -5.956695973873e-02*(V(u23_10) + V(u24_10))
+ + -1.089849546552e-01*(V(u23_11) + V(u24_11)) + -1.598252058029e-01*(V(u23_12) + V(u24_12)) + -5.745092034340e-02*(V(u23_13)
+ + V(u24_13)) + -1.558409035206e-01*(V(u23_14) + V(u24_14)) + -1.194234713912e-01*(V(u23_15) + V(u24_15))
+ + 1.153195500374e-01*(V(u23_16) + V(u24_16)) + -3.918054699898e-02*(V(u23_17) + V(u24_17)) + -1.921595633030e-01*(V(u23_18)
+ + V(u24_18)) + 1.130983531475e-01*(V(u23_19) + V(u24_19)))
B_u32_38 u32_38 0 V = tanh_psi(1.946437358856e-02 + 1.563329994678e-01*(V(u23_0) + V(u24_0)) + 2.851659059525e-02*(V(u23_1) + V(u24_1))
+ + 2.163542509079e-01*(V(u23_2) + V(u24_2)) + -1.663891971111e-02*(V(u23_3) + V(u24_3)) + 8.287215232849e-02*(V(u23_4) + V(u24_4))
+ + 1.576299965382e-01*(V(u23_5) + V(u24_5)) + 1.753807663918e-01*(V(u23_6) + V(u24_6)) + -2.075953334570e-01*(V(u23_7) + V(u24_7))
+ + 1.160400807858e-01*(V(u23_8) + V(u24_8)) + -3.056426346302e-02*(V(u23_9) + V(u24_9)) + -1.519255042076e-01*(V(u23_10) + V(u24_10))
+ + -3.484435379505e-02*(V(u23_11) + V(u24_11)) + 5.358448624611e-02*(V(u23_12) + V(u24_12)) + -1.374185085297e-01*(V(u23_13)
+ + V(u24_13)) + -6.924968957901e-02*(V(u23_14) + V(u24_14)) + 4.415124654770e-02*(V(u23_15) + V(u24_15))
+ + 1.915910840034e-01*(V(u23_16) + V(u24_16)) + -1.050768643618e-01*(V(u23_17) + V(u24_17)) + 2.119433879852e-01*(V(u23_18)
+ + V(u24_18)) + -8.586502075195e-02*(V(u23_19) + V(u24_19)))
B_u32_39 u32_39 0 V = tanh_psi(-2.926414310932e-01 + -2.042137980461e-01*(V(u23_0) + V(u24_0)) + 1.655678451061e-01*(V(u23_1) + V(u24_1))
+ + 2.182444930077e-02*(V(u23_2) + V(u24_2)) + 1.109732091427e-01*(V(u23_3) + V(u24_3)) + 2.179311215878e-01*(V(u23_4) + V(u24_4))
+ + -1.697469204664e-01*(V(u23_5) + V(u24_5)) + -4.406298696995e-02*(V(u23_6) + V(u24_6)) + 1.884983181953e-01*(V(u23_7) + V(u24_7))
+ + 2.181922793388e-01*(V(u23_8) + V(u24_8)) + -4.153238236904e-02*(V(u23_9) + V(u24_9)) + 1.289189159870e-01*(V(u23_10) + V(u24_10))
+ + -1.027061045170e-01*(V(u23_11) + V(u24_11)) + 1.858378052711e-01*(V(u23_12) + V(u24_12)) + -9.171903133392e-03*(V(u23_13)
+ + V(u24_13)) + -1.568247824907e-01*(V(u23_14) + V(u24_14)) + 1.398643553257e-01*(V(u23_15) + V(u24_15))
+ + -3.899210691452e-02*(V(u23_16) + V(u24_16)) + -1.555541753769e-01*(V(u23_17) + V(u24_17)) + 1.599707901478e-01*(V(u23_18)
+ + V(u24_18)) + -3.060330450535e-02*(V(u23_19) + V(u24_19)))
B_out_0 out0 0 V = (-8.562895655632e-02 + -1.626914739609e-02*V(u32_0) + 5.891531705856e-02*V(u32_1) + -6.724733859301e-02*V(u32_2)
+ + -1.828812062740e-02*V(u32_3) + 1.285609751940e-01*V(u32_4) + -9.111735969782e-02*V(u32_5) + -1.404555290937e-01*V(u32_6)
+ + -2.081029117107e-02*V(u32_7) + -9.755048155785e-02*V(u32_8) + 5.730369687080e-02*V(u32_9) + -1.316990405321e-01*V(u32_10)
+ + -5.221426486969e-02*V(u32_11) + -1.128220409155e-01*V(u32_12) + -5.568876862526e-02*V(u32_13) + 1.467639654875e-01*V(u32_14)
+ + -2.868589758873e-02*V(u32_15) + -1.713494956493e-02*V(u32_16) + -1.555891185999e-01*V(u32_17) + -8.687560260296e-02*V(u32_18)
+ + 1.249730139971e-01*V(u32_19) + -2.880784869194e-02*V(u32_20) + 1.190001219511e-01*V(u32_21) + 1.465555280447e-01*V(u32_22)
+ + 1.261589974165e-01*V(u32_23) + 4.593762755394e-02*V(u32_24) + -1.982197165489e-03*V(u32_25) + 6.491152942181e-02*V(u32_26)
+ + 1.876816153526e-03*V(u32_27) + -1.467765718699e-01*V(u32_28) + 1.108114868402e-01*V(u32_29) + 1.206716895103e-02*V(u32_30)
+ + -9.163775295019e-02*V(u32_31) + -2.844065427780e-03*V(u32_32) + 9.255661070347e-02*V(u32_33) + 1.291987150908e-01*V(u32_34)
+ + -4.955576360226e-02*V(u32_35) + -4.411142319441e-02*V(u32_36) + 1.010902971029e-01*V(u32_37) + -1.350494325161e-01*V(u32_38)
+ + -3.464847803116e-02*V(u32_39))

.ends psi_nn_psinn_laplace
